`default_nettype none
module life_stat(input wire clk_in,
                 input wire alive_in,
                 output logic[2*LOG_BOARD_SIZE-1:0] count_out);
endmodule
`default_nettype wire
