`default_nettype none
module life_rule(input wire[8:0] window_in,
                 output wire alive_out);
endmodule
`default_nettype wire
