module audio(input wire clk_in,
             input wire rst_in,
             input wire play_audio_in,
             output logic aud_pwm);
             

                 
 

endmodule