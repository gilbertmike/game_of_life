`include "common.svh"

`default_nettype none
module synchronizer(input wire clk_in,
                    input wire logic_done_in, render_done_in,
                    output logic logic_start_out, render_start_out,
                    output logic buf_swap_out);
endmodule
`default_nettype wire
