`timescale 1ns / 1ps

`include "common.svh"

module audio_tb(
    
    );
endmodule
