`default_nettype none
module top_level(

    );
endmodule
`default_nettype wire
