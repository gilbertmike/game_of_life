`default_nettype none
module b52bomber(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd5, 6'd18}: alive_out = 1;
            {6'd5, 6'd19}: alive_out = 1;
            {6'd5, 6'd22}: alive_out = 1;
            {6'd5, 6'd28}: alive_out = 1;
            {6'd5, 6'd29}: alive_out = 1;
            {6'd6, 6'd14}: alive_out = 1;
            {6'd6, 6'd15}: alive_out = 1;
            {6'd6, 6'd18}: alive_out = 1;
            {6'd6, 6'd19}: alive_out = 1;
            {6'd6, 6'd23}: alive_out = 1;
            {6'd6, 6'd27}: alive_out = 1;
            {6'd6, 6'd30}: alive_out = 1;
            {6'd7, 6'd14}: alive_out = 1;
            {6'd7, 6'd15}: alive_out = 1;
            {6'd7, 6'd23}: alive_out = 1;
            {6'd7, 6'd27}: alive_out = 1;
            {6'd7, 6'd29}: alive_out = 1;
            {6'd7, 6'd32}: alive_out = 1;
            {6'd8, 6'd19}: alive_out = 1;
            {6'd8, 6'd20}: alive_out = 1;
            {6'd8, 6'd21}: alive_out = 1;
            {6'd8, 6'd22}: alive_out = 1;
            {6'd8, 6'd28}: alive_out = 1;
            {6'd9, 6'd29}: alive_out = 1;
            {6'd9, 6'd30}: alive_out = 1;
            {6'd9, 6'd32}: alive_out = 1;
            {6'd10, 6'd31}: alive_out = 1;
            {6'd14, 6'd18}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd15, 6'd18}: alive_out = 1;
            {6'd15, 6'd19}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd23, 6'd31}: alive_out = 1;
            {6'd23, 6'd33}: alive_out = 1;
            {6'd24, 6'd16}: alive_out = 1;
            {6'd24, 6'd32}: alive_out = 1;
            {6'd25, 6'd15}: alive_out = 1;
            {6'd25, 6'd17}: alive_out = 1;
            {6'd26, 6'd16}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd24}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd27, 6'd31}: alive_out = 1;
            {6'd28, 6'd24}: alive_out = 1;
            {6'd28, 6'd29}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd32, 6'd20}: alive_out = 1;
            {6'd32, 6'd21}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd22}: alive_out = 1;
            {6'd33, 6'd29}: alive_out = 1;
            {6'd33, 6'd30}: alive_out = 1;
            {6'd34, 6'd29}: alive_out = 1;
            {6'd34, 6'd30}: alive_out = 1;
            {6'd38, 6'd17}: alive_out = 1;
            {6'd39, 6'd16}: alive_out = 1;
            {6'd39, 6'd18}: alive_out = 1;
            {6'd39, 6'd19}: alive_out = 1;
            {6'd40, 6'd20}: alive_out = 1;
            {6'd40, 6'd29}: alive_out = 1;
            {6'd40, 6'd30}: alive_out = 1;
            {6'd40, 6'd33}: alive_out = 1;
            {6'd41, 6'd16}: alive_out = 1;
            {6'd41, 6'd19}: alive_out = 1;
            {6'd41, 6'd21}: alive_out = 1;
            {6'd41, 6'd25}: alive_out = 1;
            {6'd41, 6'd26}: alive_out = 1;
            {6'd41, 6'd29}: alive_out = 1;
            {6'd41, 6'd30}: alive_out = 1;
            {6'd41, 6'd34}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd42, 6'd21}: alive_out = 1;
            {6'd42, 6'd25}: alive_out = 1;
            {6'd42, 6'd26}: alive_out = 1;
            {6'd42, 6'd34}: alive_out = 1;
            {6'd43, 6'd19}: alive_out = 1;
            {6'd43, 6'd20}: alive_out = 1;
            {6'd43, 6'd30}: alive_out = 1;
            {6'd43, 6'd31}: alive_out = 1;
            {6'd43, 6'd32}: alive_out = 1;
            {6'd43, 6'd33}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module shipinabottle(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd16, 6'd20}: alive_out = 1;
            {6'd16, 6'd21}: alive_out = 1;
            {6'd16, 6'd28}: alive_out = 1;
            {6'd16, 6'd29}: alive_out = 1;
            {6'd17, 6'd19}: alive_out = 1;
            {6'd17, 6'd22}: alive_out = 1;
            {6'd17, 6'd27}: alive_out = 1;
            {6'd17, 6'd30}: alive_out = 1;
            {6'd18, 6'd19}: alive_out = 1;
            {6'd18, 6'd21}: alive_out = 1;
            {6'd18, 6'd28}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd19, 6'd17}: alive_out = 1;
            {6'd19, 6'd18}: alive_out = 1;
            {6'd19, 6'd21}: alive_out = 1;
            {6'd19, 6'd22}: alive_out = 1;
            {6'd19, 6'd23}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd19, 6'd28}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd20, 6'd16}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd33}: alive_out = 1;
            {6'd21, 6'd16}: alive_out = 1;
            {6'd21, 6'd18}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd30}: alive_out = 1;
            {6'd21, 6'd31}: alive_out = 1;
            {6'd21, 6'd33}: alive_out = 1;
            {6'd22, 6'd17}: alive_out = 1;
            {6'd22, 6'd19}: alive_out = 1;
            {6'd22, 6'd30}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd23, 6'd19}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd25}: alive_out = 1;
            {6'd23, 6'd29}: alive_out = 1;
            {6'd23, 6'd30}: alive_out = 1;
            {6'd24, 6'd23}: alive_out = 1;
            {6'd24, 6'd25}: alive_out = 1;
            {6'd25, 6'd23}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd26, 6'd30}: alive_out = 1;
            {6'd27, 6'd17}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd27, 6'd32}: alive_out = 1;
            {6'd28, 6'd16}: alive_out = 1;
            {6'd28, 6'd18}: alive_out = 1;
            {6'd28, 6'd19}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd28, 6'd31}: alive_out = 1;
            {6'd28, 6'd33}: alive_out = 1;
            {6'd29, 6'd16}: alive_out = 1;
            {6'd29, 6'd23}: alive_out = 1;
            {6'd29, 6'd26}: alive_out = 1;
            {6'd29, 6'd33}: alive_out = 1;
            {6'd30, 6'd17}: alive_out = 1;
            {6'd30, 6'd18}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd30, 6'd22}: alive_out = 1;
            {6'd30, 6'd23}: alive_out = 1;
            {6'd30, 6'd26}: alive_out = 1;
            {6'd30, 6'd27}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd31}: alive_out = 1;
            {6'd30, 6'd32}: alive_out = 1;
            {6'd31, 6'd19}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd31, 6'd30}: alive_out = 1;
            {6'd32, 6'd19}: alive_out = 1;
            {6'd32, 6'd22}: alive_out = 1;
            {6'd32, 6'd27}: alive_out = 1;
            {6'd32, 6'd30}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd28}: alive_out = 1;
            {6'd33, 6'd29}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module loaflipflop(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd17}: alive_out = 1;
            {6'd9, 6'd16}: alive_out = 1;
            {6'd9, 6'd17}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd12, 6'd16}: alive_out = 1;
            {6'd12, 6'd17}: alive_out = 1;
            {6'd12, 6'd18}: alive_out = 1;
            {6'd14, 6'd16}: alive_out = 1;
            {6'd14, 6'd18}: alive_out = 1;
            {6'd15, 6'd16}: alive_out = 1;
            {6'd15, 6'd18}: alive_out = 1;
            {6'd17, 6'd16}: alive_out = 1;
            {6'd17, 6'd17}: alive_out = 1;
            {6'd17, 6'd18}: alive_out = 1;
            {6'd20, 6'd16}: alive_out = 1;
            {6'd20, 6'd17}: alive_out = 1;
            {6'd20, 6'd18}: alive_out = 1;
            {6'd21, 6'd17}: alive_out = 1;
            {6'd23, 6'd9}: alive_out = 1;
            {6'd23, 6'd10}: alive_out = 1;
            {6'd23, 6'd11}: alive_out = 1;
            {6'd23, 6'd12}: alive_out = 1;
            {6'd23, 6'd13}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd29}: alive_out = 1;
            {6'd24, 6'd8}: alive_out = 1;
            {6'd24, 6'd9}: alive_out = 1;
            {6'd24, 6'd10}: alive_out = 1;
            {6'd24, 6'd13}: alive_out = 1;
            {6'd24, 6'd14}: alive_out = 1;
            {6'd24, 6'd15}: alive_out = 1;
            {6'd24, 6'd18}: alive_out = 1;
            {6'd24, 6'd19}: alive_out = 1;
            {6'd24, 6'd27}: alive_out = 1;
            {6'd24, 6'd30}: alive_out = 1;
            {6'd25, 6'd9}: alive_out = 1;
            {6'd25, 6'd10}: alive_out = 1;
            {6'd25, 6'd11}: alive_out = 1;
            {6'd25, 6'd12}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd25, 6'd14}: alive_out = 1;
            {6'd25, 6'd17}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd26}: alive_out = 1;
            {6'd25, 6'd31}: alive_out = 1;
            {6'd26, 6'd17}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd32}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd27, 6'd32}: alive_out = 1;
            {6'd28, 6'd25}: alive_out = 1;
            {6'd28, 6'd32}: alive_out = 1;
            {6'd29, 6'd26}: alive_out = 1;
            {6'd29, 6'd31}: alive_out = 1;
            {6'd30, 6'd27}: alive_out = 1;
            {6'd30, 6'd30}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd32, 6'd19}: alive_out = 1;
            {6'd32, 6'd20}: alive_out = 1;
            {6'd32, 6'd21}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;
            {6'd33, 6'd22}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd36, 6'd16}: alive_out = 1;
            {6'd36, 6'd24}: alive_out = 1;
            {6'd37, 6'd16}: alive_out = 1;
            {6'd37, 6'd24}: alive_out = 1;
            {6'd39, 6'd17}: alive_out = 1;
            {6'd39, 6'd23}: alive_out = 1;
            {6'd40, 6'd18}: alive_out = 1;
            {6'd40, 6'd22}: alive_out = 1;
            {6'd41, 6'd19}: alive_out = 1;
            {6'd41, 6'd20}: alive_out = 1;
            {6'd41, 6'd21}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module ringoffire(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd24}: alive_out = 1;
            {6'd8, 6'd26}: alive_out = 1;
            {6'd9, 6'd22}: alive_out = 1;
            {6'd9, 6'd25}: alive_out = 1;
            {6'd9, 6'd28}: alive_out = 1;
            {6'd10, 6'd20}: alive_out = 1;
            {6'd10, 6'd23}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd10, 6'd27}: alive_out = 1;
            {6'd10, 6'd30}: alive_out = 1;
            {6'd11, 6'd18}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd11, 6'd23}: alive_out = 1;
            {6'd11, 6'd25}: alive_out = 1;
            {6'd11, 6'd27}: alive_out = 1;
            {6'd11, 6'd29}: alive_out = 1;
            {6'd11, 6'd32}: alive_out = 1;
            {6'd12, 6'd16}: alive_out = 1;
            {6'd12, 6'd19}: alive_out = 1;
            {6'd12, 6'd21}: alive_out = 1;
            {6'd12, 6'd23}: alive_out = 1;
            {6'd12, 6'd26}: alive_out = 1;
            {6'd12, 6'd29}: alive_out = 1;
            {6'd12, 6'd31}: alive_out = 1;
            {6'd13, 6'd17}: alive_out = 1;
            {6'd13, 6'd19}: alive_out = 1;
            {6'd13, 6'd22}: alive_out = 1;
            {6'd13, 6'd23}: alive_out = 1;
            {6'd13, 6'd29}: alive_out = 1;
            {6'd13, 6'd31}: alive_out = 1;
            {6'd13, 6'd32}: alive_out = 1;
            {6'd13, 6'd33}: alive_out = 1;
            {6'd14, 6'd15}: alive_out = 1;
            {6'd14, 6'd16}: alive_out = 1;
            {6'd14, 6'd17}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd30}: alive_out = 1;
            {6'd15, 6'd18}: alive_out = 1;
            {6'd15, 6'd31}: alive_out = 1;
            {6'd15, 6'd32}: alive_out = 1;
            {6'd15, 6'd33}: alive_out = 1;
            {6'd15, 6'd34}: alive_out = 1;
            {6'd16, 6'd14}: alive_out = 1;
            {6'd16, 6'd15}: alive_out = 1;
            {6'd16, 6'd16}: alive_out = 1;
            {6'd16, 6'd17}: alive_out = 1;
            {6'd17, 6'd33}: alive_out = 1;
            {6'd17, 6'd34}: alive_out = 1;
            {6'd17, 6'd35}: alive_out = 1;
            {6'd18, 6'd13}: alive_out = 1;
            {6'd18, 6'd14}: alive_out = 1;
            {6'd18, 6'd15}: alive_out = 1;
            {6'd18, 6'd32}: alive_out = 1;
            {6'd19, 6'd16}: alive_out = 1;
            {6'd19, 6'd33}: alive_out = 1;
            {6'd19, 6'd34}: alive_out = 1;
            {6'd19, 6'd35}: alive_out = 1;
            {6'd19, 6'd36}: alive_out = 1;
            {6'd20, 6'd12}: alive_out = 1;
            {6'd20, 6'd13}: alive_out = 1;
            {6'd20, 6'd14}: alive_out = 1;
            {6'd20, 6'd15}: alive_out = 1;
            {6'd21, 6'd35}: alive_out = 1;
            {6'd21, 6'd36}: alive_out = 1;
            {6'd21, 6'd37}: alive_out = 1;
            {6'd22, 6'd11}: alive_out = 1;
            {6'd22, 6'd12}: alive_out = 1;
            {6'd22, 6'd13}: alive_out = 1;
            {6'd22, 6'd34}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd23, 6'd36}: alive_out = 1;
            {6'd23, 6'd37}: alive_out = 1;
            {6'd23, 6'd38}: alive_out = 1;
            {6'd24, 6'd10}: alive_out = 1;
            {6'd24, 6'd11}: alive_out = 1;
            {6'd24, 6'd12}: alive_out = 1;
            {6'd24, 6'd13}: alive_out = 1;
            {6'd24, 6'd14}: alive_out = 1;
            {6'd25, 6'd35}: alive_out = 1;
            {6'd25, 6'd36}: alive_out = 1;
            {6'd25, 6'd37}: alive_out = 1;
            {6'd25, 6'd38}: alive_out = 1;
            {6'd25, 6'd39}: alive_out = 1;
            {6'd26, 6'd11}: alive_out = 1;
            {6'd26, 6'd12}: alive_out = 1;
            {6'd26, 6'd13}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd35}: alive_out = 1;
            {6'd27, 6'd15}: alive_out = 1;
            {6'd27, 6'd36}: alive_out = 1;
            {6'd27, 6'd37}: alive_out = 1;
            {6'd27, 6'd38}: alive_out = 1;
            {6'd28, 6'd12}: alive_out = 1;
            {6'd28, 6'd13}: alive_out = 1;
            {6'd28, 6'd14}: alive_out = 1;
            {6'd29, 6'd34}: alive_out = 1;
            {6'd29, 6'd35}: alive_out = 1;
            {6'd29, 6'd36}: alive_out = 1;
            {6'd29, 6'd37}: alive_out = 1;
            {6'd30, 6'd13}: alive_out = 1;
            {6'd30, 6'd14}: alive_out = 1;
            {6'd30, 6'd15}: alive_out = 1;
            {6'd30, 6'd16}: alive_out = 1;
            {6'd30, 6'd33}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd34}: alive_out = 1;
            {6'd31, 6'd35}: alive_out = 1;
            {6'd31, 6'd36}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd15}: alive_out = 1;
            {6'd32, 6'd16}: alive_out = 1;
            {6'd33, 6'd32}: alive_out = 1;
            {6'd33, 6'd33}: alive_out = 1;
            {6'd33, 6'd34}: alive_out = 1;
            {6'd33, 6'd35}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd16}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd35, 6'd30}: alive_out = 1;
            {6'd35, 6'd32}: alive_out = 1;
            {6'd35, 6'd33}: alive_out = 1;
            {6'd35, 6'd34}: alive_out = 1;
            {6'd36, 6'd16}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd36, 6'd26}: alive_out = 1;
            {6'd36, 6'd27}: alive_out = 1;
            {6'd36, 6'd30}: alive_out = 1;
            {6'd36, 6'd32}: alive_out = 1;
            {6'd37, 6'd18}: alive_out = 1;
            {6'd37, 6'd20}: alive_out = 1;
            {6'd37, 6'd23}: alive_out = 1;
            {6'd37, 6'd26}: alive_out = 1;
            {6'd37, 6'd28}: alive_out = 1;
            {6'd37, 6'd30}: alive_out = 1;
            {6'd37, 6'd33}: alive_out = 1;
            {6'd38, 6'd17}: alive_out = 1;
            {6'd38, 6'd20}: alive_out = 1;
            {6'd38, 6'd22}: alive_out = 1;
            {6'd38, 6'd24}: alive_out = 1;
            {6'd38, 6'd26}: alive_out = 1;
            {6'd38, 6'd28}: alive_out = 1;
            {6'd38, 6'd31}: alive_out = 1;
            {6'd39, 6'd19}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd39, 6'd24}: alive_out = 1;
            {6'd39, 6'd26}: alive_out = 1;
            {6'd39, 6'd29}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;
            {6'd40, 6'd24}: alive_out = 1;
            {6'd40, 6'd27}: alive_out = 1;
            {6'd41, 6'd23}: alive_out = 1;
            {6'd41, 6'd25}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module frothingpuffer(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd21}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd9, 6'd19}: alive_out = 1;
            {6'd9, 6'd20}: alive_out = 1;
            {6'd9, 6'd21}: alive_out = 1;
            {6'd10, 6'd18}: alive_out = 1;
            {6'd10, 6'd19}: alive_out = 1;
            {6'd10, 6'd20}: alive_out = 1;
            {6'd11, 6'd16}: alive_out = 1;
            {6'd11, 6'd20}: alive_out = 1;
            {6'd12, 6'd16}: alive_out = 1;
            {6'd12, 6'd17}: alive_out = 1;
            {6'd12, 6'd18}: alive_out = 1;
            {6'd13, 6'd15}: alive_out = 1;
            {6'd13, 6'd20}: alive_out = 1;
            {6'd13, 6'd31}: alive_out = 1;
            {6'd14, 6'd14}: alive_out = 1;
            {6'd14, 6'd15}: alive_out = 1;
            {6'd14, 6'd16}: alive_out = 1;
            {6'd14, 6'd17}: alive_out = 1;
            {6'd14, 6'd18}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd28}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd14, 6'd31}: alive_out = 1;
            {6'd15, 6'd13}: alive_out = 1;
            {6'd15, 6'd14}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd15, 6'd26}: alive_out = 1;
            {6'd15, 6'd27}: alive_out = 1;
            {6'd15, 6'd28}: alive_out = 1;
            {6'd16, 6'd14}: alive_out = 1;
            {6'd16, 6'd18}: alive_out = 1;
            {6'd16, 6'd19}: alive_out = 1;
            {6'd16, 6'd25}: alive_out = 1;
            {6'd16, 6'd26}: alive_out = 1;
            {6'd17, 6'd16}: alive_out = 1;
            {6'd17, 6'd17}: alive_out = 1;
            {6'd17, 6'd20}: alive_out = 1;
            {6'd17, 6'd23}: alive_out = 1;
            {6'd17, 6'd27}: alive_out = 1;
            {6'd17, 6'd29}: alive_out = 1;
            {6'd17, 6'd30}: alive_out = 1;
            {6'd17, 6'd32}: alive_out = 1;
            {6'd18, 6'd16}: alive_out = 1;
            {6'd18, 6'd18}: alive_out = 1;
            {6'd18, 6'd23}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd18, 6'd33}: alive_out = 1;
            {6'd19, 6'd15}: alive_out = 1;
            {6'd19, 6'd16}: alive_out = 1;
            {6'd19, 6'd17}: alive_out = 1;
            {6'd19, 6'd21}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd19, 6'd28}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd19, 6'd35}: alive_out = 1;
            {6'd20, 6'd15}: alive_out = 1;
            {6'd20, 6'd21}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd20, 6'd32}: alive_out = 1;
            {6'd20, 6'd33}: alive_out = 1;
            {6'd20, 6'd34}: alive_out = 1;
            {6'd21, 6'd15}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd27}: alive_out = 1;
            {6'd21, 6'd29}: alive_out = 1;
            {6'd21, 6'd35}: alive_out = 1;
            {6'd22, 6'd16}: alive_out = 1;
            {6'd22, 6'd20}: alive_out = 1;
            {6'd22, 6'd21}: alive_out = 1;
            {6'd22, 6'd27}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd23, 6'd17}: alive_out = 1;
            {6'd23, 6'd18}: alive_out = 1;
            {6'd23, 6'd27}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd29}: alive_out = 1;
            {6'd23, 6'd30}: alive_out = 1;
            {6'd23, 6'd31}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd21}: alive_out = 1;
            {6'd24, 6'd33}: alive_out = 1;
            {6'd25, 6'd17}: alive_out = 1;
            {6'd25, 6'd18}: alive_out = 1;
            {6'd25, 6'd27}: alive_out = 1;
            {6'd25, 6'd28}: alive_out = 1;
            {6'd25, 6'd29}: alive_out = 1;
            {6'd25, 6'd30}: alive_out = 1;
            {6'd25, 6'd31}: alive_out = 1;
            {6'd25, 6'd34}: alive_out = 1;
            {6'd26, 6'd16}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd21}: alive_out = 1;
            {6'd26, 6'd27}: alive_out = 1;
            {6'd26, 6'd32}: alive_out = 1;
            {6'd26, 6'd33}: alive_out = 1;
            {6'd27, 6'd15}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd27}: alive_out = 1;
            {6'd27, 6'd29}: alive_out = 1;
            {6'd27, 6'd35}: alive_out = 1;
            {6'd28, 6'd15}: alive_out = 1;
            {6'd28, 6'd21}: alive_out = 1;
            {6'd28, 6'd22}: alive_out = 1;
            {6'd28, 6'd23}: alive_out = 1;
            {6'd28, 6'd32}: alive_out = 1;
            {6'd28, 6'd33}: alive_out = 1;
            {6'd28, 6'd34}: alive_out = 1;
            {6'd29, 6'd15}: alive_out = 1;
            {6'd29, 6'd16}: alive_out = 1;
            {6'd29, 6'd17}: alive_out = 1;
            {6'd29, 6'd21}: alive_out = 1;
            {6'd29, 6'd27}: alive_out = 1;
            {6'd29, 6'd28}: alive_out = 1;
            {6'd29, 6'd31}: alive_out = 1;
            {6'd29, 6'd32}: alive_out = 1;
            {6'd29, 6'd35}: alive_out = 1;
            {6'd30, 6'd16}: alive_out = 1;
            {6'd30, 6'd18}: alive_out = 1;
            {6'd30, 6'd23}: alive_out = 1;
            {6'd30, 6'd24}: alive_out = 1;
            {6'd30, 6'd25}: alive_out = 1;
            {6'd30, 6'd30}: alive_out = 1;
            {6'd30, 6'd33}: alive_out = 1;
            {6'd31, 6'd16}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd20}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd31, 6'd27}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd31, 6'd30}: alive_out = 1;
            {6'd31, 6'd32}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd18}: alive_out = 1;
            {6'd32, 6'd19}: alive_out = 1;
            {6'd32, 6'd25}: alive_out = 1;
            {6'd32, 6'd26}: alive_out = 1;
            {6'd33, 6'd13}: alive_out = 1;
            {6'd33, 6'd14}: alive_out = 1;
            {6'd33, 6'd25}: alive_out = 1;
            {6'd33, 6'd26}: alive_out = 1;
            {6'd33, 6'd27}: alive_out = 1;
            {6'd33, 6'd28}: alive_out = 1;
            {6'd34, 6'd14}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd16}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd19}: alive_out = 1;
            {6'd34, 6'd28}: alive_out = 1;
            {6'd34, 6'd29}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd35, 6'd15}: alive_out = 1;
            {6'd35, 6'd20}: alive_out = 1;
            {6'd35, 6'd31}: alive_out = 1;
            {6'd36, 6'd16}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd37, 6'd16}: alive_out = 1;
            {6'd37, 6'd20}: alive_out = 1;
            {6'd38, 6'd18}: alive_out = 1;
            {6'd38, 6'd19}: alive_out = 1;
            {6'd38, 6'd20}: alive_out = 1;
            {6'd39, 6'd18}: alive_out = 1;
            {6'd39, 6'd19}: alive_out = 1;
            {6'd39, 6'd20}: alive_out = 1;
            {6'd39, 6'd21}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module venetial_blinds(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd6, 6'd2}: alive_out = 1;
            {6'd6, 6'd3}: alive_out = 1;
            {6'd6, 6'd4}: alive_out = 1;
            {6'd6, 6'd5}: alive_out = 1;
            {6'd6, 6'd6}: alive_out = 1;
            {6'd6, 6'd7}: alive_out = 1;
            {6'd6, 6'd8}: alive_out = 1;
            {6'd6, 6'd9}: alive_out = 1;
            {6'd6, 6'd10}: alive_out = 1;
            {6'd6, 6'd11}: alive_out = 1;
            {6'd6, 6'd12}: alive_out = 1;
            {6'd6, 6'd13}: alive_out = 1;
            {6'd6, 6'd14}: alive_out = 1;
            {6'd6, 6'd15}: alive_out = 1;
            {6'd6, 6'd16}: alive_out = 1;
            {6'd6, 6'd17}: alive_out = 1;
            {6'd6, 6'd18}: alive_out = 1;
            {6'd6, 6'd19}: alive_out = 1;
            {6'd6, 6'd20}: alive_out = 1;
            {6'd6, 6'd21}: alive_out = 1;
            {6'd6, 6'd22}: alive_out = 1;
            {6'd6, 6'd23}: alive_out = 1;
            {6'd6, 6'd24}: alive_out = 1;
            {6'd6, 6'd25}: alive_out = 1;
            {6'd6, 6'd26}: alive_out = 1;
            {6'd6, 6'd27}: alive_out = 1;
            {6'd6, 6'd28}: alive_out = 1;
            {6'd6, 6'd29}: alive_out = 1;
            {6'd6, 6'd30}: alive_out = 1;
            {6'd6, 6'd31}: alive_out = 1;
            {6'd6, 6'd32}: alive_out = 1;
            {6'd6, 6'd33}: alive_out = 1;
            {6'd6, 6'd34}: alive_out = 1;
            {6'd6, 6'd35}: alive_out = 1;
            {6'd6, 6'd36}: alive_out = 1;
            {6'd6, 6'd37}: alive_out = 1;
            {6'd6, 6'd38}: alive_out = 1;
            {6'd6, 6'd39}: alive_out = 1;
            {6'd6, 6'd40}: alive_out = 1;
            {6'd6, 6'd41}: alive_out = 1;
            {6'd6, 6'd42}: alive_out = 1;
            {6'd6, 6'd43}: alive_out = 1;
            {6'd6, 6'd44}: alive_out = 1;
            {6'd6, 6'd45}: alive_out = 1;
            {6'd6, 6'd46}: alive_out = 1;
            {6'd7, 6'd2}: alive_out = 1;
            {6'd7, 6'd3}: alive_out = 1;
            {6'd7, 6'd4}: alive_out = 1;
            {6'd7, 6'd5}: alive_out = 1;
            {6'd7, 6'd6}: alive_out = 1;
            {6'd7, 6'd7}: alive_out = 1;
            {6'd7, 6'd8}: alive_out = 1;
            {6'd7, 6'd9}: alive_out = 1;
            {6'd7, 6'd10}: alive_out = 1;
            {6'd7, 6'd11}: alive_out = 1;
            {6'd7, 6'd12}: alive_out = 1;
            {6'd7, 6'd13}: alive_out = 1;
            {6'd7, 6'd14}: alive_out = 1;
            {6'd7, 6'd15}: alive_out = 1;
            {6'd7, 6'd16}: alive_out = 1;
            {6'd7, 6'd17}: alive_out = 1;
            {6'd7, 6'd18}: alive_out = 1;
            {6'd7, 6'd19}: alive_out = 1;
            {6'd7, 6'd20}: alive_out = 1;
            {6'd7, 6'd21}: alive_out = 1;
            {6'd7, 6'd22}: alive_out = 1;
            {6'd7, 6'd23}: alive_out = 1;
            {6'd7, 6'd24}: alive_out = 1;
            {6'd7, 6'd25}: alive_out = 1;
            {6'd7, 6'd26}: alive_out = 1;
            {6'd7, 6'd27}: alive_out = 1;
            {6'd7, 6'd28}: alive_out = 1;
            {6'd7, 6'd29}: alive_out = 1;
            {6'd7, 6'd30}: alive_out = 1;
            {6'd7, 6'd31}: alive_out = 1;
            {6'd7, 6'd32}: alive_out = 1;
            {6'd7, 6'd33}: alive_out = 1;
            {6'd7, 6'd34}: alive_out = 1;
            {6'd7, 6'd35}: alive_out = 1;
            {6'd7, 6'd36}: alive_out = 1;
            {6'd7, 6'd37}: alive_out = 1;
            {6'd7, 6'd38}: alive_out = 1;
            {6'd7, 6'd39}: alive_out = 1;
            {6'd7, 6'd40}: alive_out = 1;
            {6'd7, 6'd41}: alive_out = 1;
            {6'd7, 6'd42}: alive_out = 1;
            {6'd7, 6'd43}: alive_out = 1;
            {6'd7, 6'd44}: alive_out = 1;
            {6'd7, 6'd45}: alive_out = 1;
            {6'd7, 6'd46}: alive_out = 1;
            {6'd10, 6'd2}: alive_out = 1;
            {6'd10, 6'd3}: alive_out = 1;
            {6'd10, 6'd4}: alive_out = 1;
            {6'd10, 6'd5}: alive_out = 1;
            {6'd10, 6'd6}: alive_out = 1;
            {6'd10, 6'd7}: alive_out = 1;
            {6'd10, 6'd8}: alive_out = 1;
            {6'd10, 6'd9}: alive_out = 1;
            {6'd10, 6'd10}: alive_out = 1;
            {6'd10, 6'd11}: alive_out = 1;
            {6'd10, 6'd12}: alive_out = 1;
            {6'd10, 6'd13}: alive_out = 1;
            {6'd10, 6'd14}: alive_out = 1;
            {6'd10, 6'd15}: alive_out = 1;
            {6'd10, 6'd16}: alive_out = 1;
            {6'd10, 6'd17}: alive_out = 1;
            {6'd10, 6'd18}: alive_out = 1;
            {6'd10, 6'd19}: alive_out = 1;
            {6'd10, 6'd20}: alive_out = 1;
            {6'd10, 6'd21}: alive_out = 1;
            {6'd10, 6'd22}: alive_out = 1;
            {6'd10, 6'd23}: alive_out = 1;
            {6'd10, 6'd24}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd10, 6'd26}: alive_out = 1;
            {6'd10, 6'd27}: alive_out = 1;
            {6'd10, 6'd28}: alive_out = 1;
            {6'd10, 6'd29}: alive_out = 1;
            {6'd10, 6'd30}: alive_out = 1;
            {6'd10, 6'd31}: alive_out = 1;
            {6'd10, 6'd32}: alive_out = 1;
            {6'd10, 6'd33}: alive_out = 1;
            {6'd10, 6'd34}: alive_out = 1;
            {6'd10, 6'd35}: alive_out = 1;
            {6'd10, 6'd36}: alive_out = 1;
            {6'd10, 6'd37}: alive_out = 1;
            {6'd10, 6'd38}: alive_out = 1;
            {6'd10, 6'd39}: alive_out = 1;
            {6'd10, 6'd40}: alive_out = 1;
            {6'd10, 6'd41}: alive_out = 1;
            {6'd10, 6'd42}: alive_out = 1;
            {6'd10, 6'd43}: alive_out = 1;
            {6'd10, 6'd44}: alive_out = 1;
            {6'd10, 6'd45}: alive_out = 1;
            {6'd10, 6'd46}: alive_out = 1;
            {6'd11, 6'd2}: alive_out = 1;
            {6'd11, 6'd3}: alive_out = 1;
            {6'd11, 6'd4}: alive_out = 1;
            {6'd11, 6'd5}: alive_out = 1;
            {6'd11, 6'd6}: alive_out = 1;
            {6'd11, 6'd7}: alive_out = 1;
            {6'd11, 6'd8}: alive_out = 1;
            {6'd11, 6'd9}: alive_out = 1;
            {6'd11, 6'd10}: alive_out = 1;
            {6'd11, 6'd11}: alive_out = 1;
            {6'd11, 6'd12}: alive_out = 1;
            {6'd11, 6'd13}: alive_out = 1;
            {6'd11, 6'd14}: alive_out = 1;
            {6'd11, 6'd15}: alive_out = 1;
            {6'd11, 6'd16}: alive_out = 1;
            {6'd11, 6'd17}: alive_out = 1;
            {6'd11, 6'd18}: alive_out = 1;
            {6'd11, 6'd19}: alive_out = 1;
            {6'd11, 6'd20}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd11, 6'd22}: alive_out = 1;
            {6'd11, 6'd23}: alive_out = 1;
            {6'd11, 6'd24}: alive_out = 1;
            {6'd11, 6'd25}: alive_out = 1;
            {6'd11, 6'd26}: alive_out = 1;
            {6'd11, 6'd27}: alive_out = 1;
            {6'd11, 6'd28}: alive_out = 1;
            {6'd11, 6'd29}: alive_out = 1;
            {6'd11, 6'd30}: alive_out = 1;
            {6'd11, 6'd31}: alive_out = 1;
            {6'd11, 6'd32}: alive_out = 1;
            {6'd11, 6'd33}: alive_out = 1;
            {6'd11, 6'd34}: alive_out = 1;
            {6'd11, 6'd35}: alive_out = 1;
            {6'd11, 6'd36}: alive_out = 1;
            {6'd11, 6'd37}: alive_out = 1;
            {6'd11, 6'd38}: alive_out = 1;
            {6'd11, 6'd39}: alive_out = 1;
            {6'd11, 6'd40}: alive_out = 1;
            {6'd11, 6'd41}: alive_out = 1;
            {6'd11, 6'd42}: alive_out = 1;
            {6'd11, 6'd43}: alive_out = 1;
            {6'd11, 6'd44}: alive_out = 1;
            {6'd11, 6'd45}: alive_out = 1;
            {6'd11, 6'd46}: alive_out = 1;
            {6'd14, 6'd2}: alive_out = 1;
            {6'd14, 6'd3}: alive_out = 1;
            {6'd14, 6'd4}: alive_out = 1;
            {6'd14, 6'd5}: alive_out = 1;
            {6'd14, 6'd6}: alive_out = 1;
            {6'd14, 6'd7}: alive_out = 1;
            {6'd14, 6'd8}: alive_out = 1;
            {6'd14, 6'd9}: alive_out = 1;
            {6'd14, 6'd10}: alive_out = 1;
            {6'd14, 6'd11}: alive_out = 1;
            {6'd14, 6'd12}: alive_out = 1;
            {6'd14, 6'd13}: alive_out = 1;
            {6'd14, 6'd14}: alive_out = 1;
            {6'd14, 6'd15}: alive_out = 1;
            {6'd14, 6'd16}: alive_out = 1;
            {6'd14, 6'd17}: alive_out = 1;
            {6'd14, 6'd18}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd20}: alive_out = 1;
            {6'd14, 6'd21}: alive_out = 1;
            {6'd14, 6'd22}: alive_out = 1;
            {6'd14, 6'd23}: alive_out = 1;
            {6'd14, 6'd24}: alive_out = 1;
            {6'd14, 6'd25}: alive_out = 1;
            {6'd14, 6'd26}: alive_out = 1;
            {6'd14, 6'd27}: alive_out = 1;
            {6'd14, 6'd28}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd14, 6'd30}: alive_out = 1;
            {6'd14, 6'd31}: alive_out = 1;
            {6'd14, 6'd32}: alive_out = 1;
            {6'd14, 6'd33}: alive_out = 1;
            {6'd14, 6'd34}: alive_out = 1;
            {6'd14, 6'd35}: alive_out = 1;
            {6'd14, 6'd36}: alive_out = 1;
            {6'd14, 6'd37}: alive_out = 1;
            {6'd14, 6'd38}: alive_out = 1;
            {6'd14, 6'd39}: alive_out = 1;
            {6'd14, 6'd40}: alive_out = 1;
            {6'd14, 6'd41}: alive_out = 1;
            {6'd14, 6'd42}: alive_out = 1;
            {6'd14, 6'd43}: alive_out = 1;
            {6'd14, 6'd44}: alive_out = 1;
            {6'd14, 6'd45}: alive_out = 1;
            {6'd14, 6'd46}: alive_out = 1;
            {6'd15, 6'd2}: alive_out = 1;
            {6'd15, 6'd3}: alive_out = 1;
            {6'd15, 6'd4}: alive_out = 1;
            {6'd15, 6'd5}: alive_out = 1;
            {6'd15, 6'd6}: alive_out = 1;
            {6'd15, 6'd7}: alive_out = 1;
            {6'd15, 6'd8}: alive_out = 1;
            {6'd15, 6'd9}: alive_out = 1;
            {6'd15, 6'd10}: alive_out = 1;
            {6'd15, 6'd11}: alive_out = 1;
            {6'd15, 6'd12}: alive_out = 1;
            {6'd15, 6'd13}: alive_out = 1;
            {6'd15, 6'd14}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd15, 6'd16}: alive_out = 1;
            {6'd15, 6'd17}: alive_out = 1;
            {6'd15, 6'd18}: alive_out = 1;
            {6'd15, 6'd19}: alive_out = 1;
            {6'd15, 6'd20}: alive_out = 1;
            {6'd15, 6'd21}: alive_out = 1;
            {6'd15, 6'd22}: alive_out = 1;
            {6'd15, 6'd23}: alive_out = 1;
            {6'd15, 6'd24}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd15, 6'd26}: alive_out = 1;
            {6'd15, 6'd27}: alive_out = 1;
            {6'd15, 6'd28}: alive_out = 1;
            {6'd15, 6'd29}: alive_out = 1;
            {6'd15, 6'd30}: alive_out = 1;
            {6'd15, 6'd31}: alive_out = 1;
            {6'd15, 6'd32}: alive_out = 1;
            {6'd15, 6'd33}: alive_out = 1;
            {6'd15, 6'd34}: alive_out = 1;
            {6'd15, 6'd35}: alive_out = 1;
            {6'd15, 6'd36}: alive_out = 1;
            {6'd15, 6'd37}: alive_out = 1;
            {6'd15, 6'd38}: alive_out = 1;
            {6'd15, 6'd39}: alive_out = 1;
            {6'd15, 6'd40}: alive_out = 1;
            {6'd15, 6'd41}: alive_out = 1;
            {6'd15, 6'd42}: alive_out = 1;
            {6'd15, 6'd43}: alive_out = 1;
            {6'd15, 6'd44}: alive_out = 1;
            {6'd15, 6'd45}: alive_out = 1;
            {6'd15, 6'd46}: alive_out = 1;
            {6'd18, 6'd2}: alive_out = 1;
            {6'd18, 6'd3}: alive_out = 1;
            {6'd18, 6'd4}: alive_out = 1;
            {6'd18, 6'd5}: alive_out = 1;
            {6'd18, 6'd6}: alive_out = 1;
            {6'd18, 6'd7}: alive_out = 1;
            {6'd18, 6'd8}: alive_out = 1;
            {6'd18, 6'd9}: alive_out = 1;
            {6'd18, 6'd10}: alive_out = 1;
            {6'd18, 6'd11}: alive_out = 1;
            {6'd18, 6'd12}: alive_out = 1;
            {6'd18, 6'd13}: alive_out = 1;
            {6'd18, 6'd14}: alive_out = 1;
            {6'd18, 6'd15}: alive_out = 1;
            {6'd18, 6'd16}: alive_out = 1;
            {6'd18, 6'd17}: alive_out = 1;
            {6'd18, 6'd18}: alive_out = 1;
            {6'd18, 6'd19}: alive_out = 1;
            {6'd18, 6'd20}: alive_out = 1;
            {6'd18, 6'd21}: alive_out = 1;
            {6'd18, 6'd22}: alive_out = 1;
            {6'd18, 6'd23}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd18, 6'd26}: alive_out = 1;
            {6'd18, 6'd27}: alive_out = 1;
            {6'd18, 6'd28}: alive_out = 1;
            {6'd18, 6'd29}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd18, 6'd31}: alive_out = 1;
            {6'd18, 6'd32}: alive_out = 1;
            {6'd18, 6'd33}: alive_out = 1;
            {6'd18, 6'd34}: alive_out = 1;
            {6'd18, 6'd35}: alive_out = 1;
            {6'd18, 6'd36}: alive_out = 1;
            {6'd18, 6'd37}: alive_out = 1;
            {6'd18, 6'd38}: alive_out = 1;
            {6'd18, 6'd39}: alive_out = 1;
            {6'd18, 6'd40}: alive_out = 1;
            {6'd18, 6'd41}: alive_out = 1;
            {6'd18, 6'd42}: alive_out = 1;
            {6'd18, 6'd43}: alive_out = 1;
            {6'd18, 6'd44}: alive_out = 1;
            {6'd18, 6'd45}: alive_out = 1;
            {6'd18, 6'd46}: alive_out = 1;
            {6'd19, 6'd2}: alive_out = 1;
            {6'd19, 6'd3}: alive_out = 1;
            {6'd19, 6'd4}: alive_out = 1;
            {6'd19, 6'd5}: alive_out = 1;
            {6'd19, 6'd6}: alive_out = 1;
            {6'd19, 6'd7}: alive_out = 1;
            {6'd19, 6'd8}: alive_out = 1;
            {6'd19, 6'd9}: alive_out = 1;
            {6'd19, 6'd10}: alive_out = 1;
            {6'd19, 6'd11}: alive_out = 1;
            {6'd19, 6'd12}: alive_out = 1;
            {6'd19, 6'd13}: alive_out = 1;
            {6'd19, 6'd14}: alive_out = 1;
            {6'd19, 6'd15}: alive_out = 1;
            {6'd19, 6'd16}: alive_out = 1;
            {6'd19, 6'd17}: alive_out = 1;
            {6'd19, 6'd18}: alive_out = 1;
            {6'd19, 6'd19}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd19, 6'd21}: alive_out = 1;
            {6'd19, 6'd22}: alive_out = 1;
            {6'd19, 6'd23}: alive_out = 1;
            {6'd19, 6'd24}: alive_out = 1;
            {6'd19, 6'd25}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd19, 6'd28}: alive_out = 1;
            {6'd19, 6'd29}: alive_out = 1;
            {6'd19, 6'd30}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd19, 6'd33}: alive_out = 1;
            {6'd19, 6'd34}: alive_out = 1;
            {6'd19, 6'd35}: alive_out = 1;
            {6'd19, 6'd36}: alive_out = 1;
            {6'd19, 6'd37}: alive_out = 1;
            {6'd19, 6'd38}: alive_out = 1;
            {6'd19, 6'd39}: alive_out = 1;
            {6'd19, 6'd40}: alive_out = 1;
            {6'd19, 6'd41}: alive_out = 1;
            {6'd19, 6'd42}: alive_out = 1;
            {6'd19, 6'd43}: alive_out = 1;
            {6'd19, 6'd44}: alive_out = 1;
            {6'd19, 6'd45}: alive_out = 1;
            {6'd19, 6'd46}: alive_out = 1;
            {6'd22, 6'd2}: alive_out = 1;
            {6'd22, 6'd3}: alive_out = 1;
            {6'd22, 6'd4}: alive_out = 1;
            {6'd22, 6'd5}: alive_out = 1;
            {6'd22, 6'd6}: alive_out = 1;
            {6'd22, 6'd7}: alive_out = 1;
            {6'd22, 6'd8}: alive_out = 1;
            {6'd22, 6'd9}: alive_out = 1;
            {6'd22, 6'd10}: alive_out = 1;
            {6'd22, 6'd11}: alive_out = 1;
            {6'd22, 6'd12}: alive_out = 1;
            {6'd22, 6'd13}: alive_out = 1;
            {6'd22, 6'd14}: alive_out = 1;
            {6'd22, 6'd15}: alive_out = 1;
            {6'd22, 6'd16}: alive_out = 1;
            {6'd22, 6'd17}: alive_out = 1;
            {6'd22, 6'd18}: alive_out = 1;
            {6'd22, 6'd19}: alive_out = 1;
            {6'd22, 6'd20}: alive_out = 1;
            {6'd22, 6'd21}: alive_out = 1;
            {6'd22, 6'd22}: alive_out = 1;
            {6'd22, 6'd23}: alive_out = 1;
            {6'd22, 6'd24}: alive_out = 1;
            {6'd22, 6'd25}: alive_out = 1;
            {6'd22, 6'd26}: alive_out = 1;
            {6'd22, 6'd27}: alive_out = 1;
            {6'd22, 6'd28}: alive_out = 1;
            {6'd22, 6'd29}: alive_out = 1;
            {6'd22, 6'd30}: alive_out = 1;
            {6'd22, 6'd31}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd22, 6'd34}: alive_out = 1;
            {6'd22, 6'd35}: alive_out = 1;
            {6'd22, 6'd36}: alive_out = 1;
            {6'd22, 6'd37}: alive_out = 1;
            {6'd22, 6'd38}: alive_out = 1;
            {6'd22, 6'd39}: alive_out = 1;
            {6'd22, 6'd40}: alive_out = 1;
            {6'd22, 6'd41}: alive_out = 1;
            {6'd22, 6'd42}: alive_out = 1;
            {6'd22, 6'd43}: alive_out = 1;
            {6'd22, 6'd44}: alive_out = 1;
            {6'd22, 6'd45}: alive_out = 1;
            {6'd22, 6'd46}: alive_out = 1;
            {6'd23, 6'd2}: alive_out = 1;
            {6'd23, 6'd3}: alive_out = 1;
            {6'd23, 6'd4}: alive_out = 1;
            {6'd23, 6'd5}: alive_out = 1;
            {6'd23, 6'd6}: alive_out = 1;
            {6'd23, 6'd7}: alive_out = 1;
            {6'd23, 6'd8}: alive_out = 1;
            {6'd23, 6'd9}: alive_out = 1;
            {6'd23, 6'd10}: alive_out = 1;
            {6'd23, 6'd11}: alive_out = 1;
            {6'd23, 6'd12}: alive_out = 1;
            {6'd23, 6'd13}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd15}: alive_out = 1;
            {6'd23, 6'd16}: alive_out = 1;
            {6'd23, 6'd17}: alive_out = 1;
            {6'd23, 6'd18}: alive_out = 1;
            {6'd23, 6'd19}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd21}: alive_out = 1;
            {6'd23, 6'd22}: alive_out = 1;
            {6'd23, 6'd23}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd25}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd23, 6'd27}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd29}: alive_out = 1;
            {6'd23, 6'd30}: alive_out = 1;
            {6'd23, 6'd31}: alive_out = 1;
            {6'd23, 6'd32}: alive_out = 1;
            {6'd23, 6'd33}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd23, 6'd36}: alive_out = 1;
            {6'd23, 6'd37}: alive_out = 1;
            {6'd23, 6'd38}: alive_out = 1;
            {6'd23, 6'd39}: alive_out = 1;
            {6'd23, 6'd40}: alive_out = 1;
            {6'd23, 6'd41}: alive_out = 1;
            {6'd23, 6'd42}: alive_out = 1;
            {6'd23, 6'd43}: alive_out = 1;
            {6'd23, 6'd44}: alive_out = 1;
            {6'd23, 6'd45}: alive_out = 1;
            {6'd23, 6'd46}: alive_out = 1;
            {6'd26, 6'd2}: alive_out = 1;
            {6'd26, 6'd3}: alive_out = 1;
            {6'd26, 6'd4}: alive_out = 1;
            {6'd26, 6'd5}: alive_out = 1;
            {6'd26, 6'd6}: alive_out = 1;
            {6'd26, 6'd7}: alive_out = 1;
            {6'd26, 6'd8}: alive_out = 1;
            {6'd26, 6'd9}: alive_out = 1;
            {6'd26, 6'd10}: alive_out = 1;
            {6'd26, 6'd11}: alive_out = 1;
            {6'd26, 6'd12}: alive_out = 1;
            {6'd26, 6'd13}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd15}: alive_out = 1;
            {6'd26, 6'd16}: alive_out = 1;
            {6'd26, 6'd17}: alive_out = 1;
            {6'd26, 6'd18}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd21}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd26}: alive_out = 1;
            {6'd26, 6'd27}: alive_out = 1;
            {6'd26, 6'd28}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd26, 6'd30}: alive_out = 1;
            {6'd26, 6'd31}: alive_out = 1;
            {6'd26, 6'd32}: alive_out = 1;
            {6'd26, 6'd33}: alive_out = 1;
            {6'd26, 6'd34}: alive_out = 1;
            {6'd26, 6'd35}: alive_out = 1;
            {6'd26, 6'd36}: alive_out = 1;
            {6'd26, 6'd37}: alive_out = 1;
            {6'd26, 6'd38}: alive_out = 1;
            {6'd26, 6'd39}: alive_out = 1;
            {6'd26, 6'd40}: alive_out = 1;
            {6'd26, 6'd41}: alive_out = 1;
            {6'd26, 6'd42}: alive_out = 1;
            {6'd26, 6'd43}: alive_out = 1;
            {6'd26, 6'd44}: alive_out = 1;
            {6'd26, 6'd45}: alive_out = 1;
            {6'd26, 6'd46}: alive_out = 1;
            {6'd27, 6'd2}: alive_out = 1;
            {6'd27, 6'd3}: alive_out = 1;
            {6'd27, 6'd4}: alive_out = 1;
            {6'd27, 6'd5}: alive_out = 1;
            {6'd27, 6'd6}: alive_out = 1;
            {6'd27, 6'd7}: alive_out = 1;
            {6'd27, 6'd8}: alive_out = 1;
            {6'd27, 6'd9}: alive_out = 1;
            {6'd27, 6'd10}: alive_out = 1;
            {6'd27, 6'd11}: alive_out = 1;
            {6'd27, 6'd12}: alive_out = 1;
            {6'd27, 6'd13}: alive_out = 1;
            {6'd27, 6'd14}: alive_out = 1;
            {6'd27, 6'd15}: alive_out = 1;
            {6'd27, 6'd16}: alive_out = 1;
            {6'd27, 6'd17}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd20}: alive_out = 1;
            {6'd27, 6'd21}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd23}: alive_out = 1;
            {6'd27, 6'd24}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd27, 6'd26}: alive_out = 1;
            {6'd27, 6'd27}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd27, 6'd29}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd27, 6'd31}: alive_out = 1;
            {6'd27, 6'd32}: alive_out = 1;
            {6'd27, 6'd33}: alive_out = 1;
            {6'd27, 6'd34}: alive_out = 1;
            {6'd27, 6'd35}: alive_out = 1;
            {6'd27, 6'd36}: alive_out = 1;
            {6'd27, 6'd37}: alive_out = 1;
            {6'd27, 6'd38}: alive_out = 1;
            {6'd27, 6'd39}: alive_out = 1;
            {6'd27, 6'd40}: alive_out = 1;
            {6'd27, 6'd41}: alive_out = 1;
            {6'd27, 6'd42}: alive_out = 1;
            {6'd27, 6'd43}: alive_out = 1;
            {6'd27, 6'd44}: alive_out = 1;
            {6'd27, 6'd45}: alive_out = 1;
            {6'd27, 6'd46}: alive_out = 1;
            {6'd30, 6'd2}: alive_out = 1;
            {6'd30, 6'd3}: alive_out = 1;
            {6'd30, 6'd4}: alive_out = 1;
            {6'd30, 6'd5}: alive_out = 1;
            {6'd30, 6'd6}: alive_out = 1;
            {6'd30, 6'd7}: alive_out = 1;
            {6'd30, 6'd8}: alive_out = 1;
            {6'd30, 6'd9}: alive_out = 1;
            {6'd30, 6'd10}: alive_out = 1;
            {6'd30, 6'd11}: alive_out = 1;
            {6'd30, 6'd12}: alive_out = 1;
            {6'd30, 6'd13}: alive_out = 1;
            {6'd30, 6'd14}: alive_out = 1;
            {6'd30, 6'd15}: alive_out = 1;
            {6'd30, 6'd16}: alive_out = 1;
            {6'd30, 6'd17}: alive_out = 1;
            {6'd30, 6'd18}: alive_out = 1;
            {6'd30, 6'd19}: alive_out = 1;
            {6'd30, 6'd20}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd30, 6'd22}: alive_out = 1;
            {6'd30, 6'd23}: alive_out = 1;
            {6'd30, 6'd24}: alive_out = 1;
            {6'd30, 6'd25}: alive_out = 1;
            {6'd30, 6'd26}: alive_out = 1;
            {6'd30, 6'd27}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd29}: alive_out = 1;
            {6'd30, 6'd30}: alive_out = 1;
            {6'd30, 6'd31}: alive_out = 1;
            {6'd30, 6'd32}: alive_out = 1;
            {6'd30, 6'd33}: alive_out = 1;
            {6'd30, 6'd34}: alive_out = 1;
            {6'd30, 6'd35}: alive_out = 1;
            {6'd30, 6'd36}: alive_out = 1;
            {6'd30, 6'd37}: alive_out = 1;
            {6'd30, 6'd38}: alive_out = 1;
            {6'd30, 6'd39}: alive_out = 1;
            {6'd30, 6'd40}: alive_out = 1;
            {6'd30, 6'd41}: alive_out = 1;
            {6'd30, 6'd42}: alive_out = 1;
            {6'd30, 6'd43}: alive_out = 1;
            {6'd30, 6'd44}: alive_out = 1;
            {6'd30, 6'd45}: alive_out = 1;
            {6'd30, 6'd46}: alive_out = 1;
            {6'd31, 6'd2}: alive_out = 1;
            {6'd31, 6'd3}: alive_out = 1;
            {6'd31, 6'd4}: alive_out = 1;
            {6'd31, 6'd5}: alive_out = 1;
            {6'd31, 6'd6}: alive_out = 1;
            {6'd31, 6'd7}: alive_out = 1;
            {6'd31, 6'd8}: alive_out = 1;
            {6'd31, 6'd9}: alive_out = 1;
            {6'd31, 6'd10}: alive_out = 1;
            {6'd31, 6'd11}: alive_out = 1;
            {6'd31, 6'd12}: alive_out = 1;
            {6'd31, 6'd13}: alive_out = 1;
            {6'd31, 6'd14}: alive_out = 1;
            {6'd31, 6'd15}: alive_out = 1;
            {6'd31, 6'd16}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd18}: alive_out = 1;
            {6'd31, 6'd19}: alive_out = 1;
            {6'd31, 6'd20}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd22}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd31, 6'd24}: alive_out = 1;
            {6'd31, 6'd25}: alive_out = 1;
            {6'd31, 6'd26}: alive_out = 1;
            {6'd31, 6'd27}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd31, 6'd30}: alive_out = 1;
            {6'd31, 6'd31}: alive_out = 1;
            {6'd31, 6'd32}: alive_out = 1;
            {6'd31, 6'd33}: alive_out = 1;
            {6'd31, 6'd34}: alive_out = 1;
            {6'd31, 6'd35}: alive_out = 1;
            {6'd31, 6'd36}: alive_out = 1;
            {6'd31, 6'd37}: alive_out = 1;
            {6'd31, 6'd38}: alive_out = 1;
            {6'd31, 6'd39}: alive_out = 1;
            {6'd31, 6'd40}: alive_out = 1;
            {6'd31, 6'd41}: alive_out = 1;
            {6'd31, 6'd42}: alive_out = 1;
            {6'd31, 6'd43}: alive_out = 1;
            {6'd31, 6'd44}: alive_out = 1;
            {6'd31, 6'd45}: alive_out = 1;
            {6'd31, 6'd46}: alive_out = 1;
            {6'd34, 6'd2}: alive_out = 1;
            {6'd34, 6'd3}: alive_out = 1;
            {6'd34, 6'd4}: alive_out = 1;
            {6'd34, 6'd5}: alive_out = 1;
            {6'd34, 6'd6}: alive_out = 1;
            {6'd34, 6'd7}: alive_out = 1;
            {6'd34, 6'd8}: alive_out = 1;
            {6'd34, 6'd9}: alive_out = 1;
            {6'd34, 6'd10}: alive_out = 1;
            {6'd34, 6'd11}: alive_out = 1;
            {6'd34, 6'd12}: alive_out = 1;
            {6'd34, 6'd13}: alive_out = 1;
            {6'd34, 6'd14}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd16}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd19}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd34, 6'd21}: alive_out = 1;
            {6'd34, 6'd22}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd34, 6'd24}: alive_out = 1;
            {6'd34, 6'd25}: alive_out = 1;
            {6'd34, 6'd26}: alive_out = 1;
            {6'd34, 6'd27}: alive_out = 1;
            {6'd34, 6'd28}: alive_out = 1;
            {6'd34, 6'd29}: alive_out = 1;
            {6'd34, 6'd30}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd34, 6'd32}: alive_out = 1;
            {6'd34, 6'd33}: alive_out = 1;
            {6'd34, 6'd34}: alive_out = 1;
            {6'd34, 6'd35}: alive_out = 1;
            {6'd34, 6'd36}: alive_out = 1;
            {6'd34, 6'd37}: alive_out = 1;
            {6'd34, 6'd38}: alive_out = 1;
            {6'd34, 6'd39}: alive_out = 1;
            {6'd34, 6'd40}: alive_out = 1;
            {6'd34, 6'd41}: alive_out = 1;
            {6'd34, 6'd42}: alive_out = 1;
            {6'd34, 6'd43}: alive_out = 1;
            {6'd34, 6'd44}: alive_out = 1;
            {6'd34, 6'd45}: alive_out = 1;
            {6'd34, 6'd46}: alive_out = 1;
            {6'd35, 6'd2}: alive_out = 1;
            {6'd35, 6'd3}: alive_out = 1;
            {6'd35, 6'd4}: alive_out = 1;
            {6'd35, 6'd5}: alive_out = 1;
            {6'd35, 6'd6}: alive_out = 1;
            {6'd35, 6'd7}: alive_out = 1;
            {6'd35, 6'd8}: alive_out = 1;
            {6'd35, 6'd9}: alive_out = 1;
            {6'd35, 6'd10}: alive_out = 1;
            {6'd35, 6'd11}: alive_out = 1;
            {6'd35, 6'd12}: alive_out = 1;
            {6'd35, 6'd13}: alive_out = 1;
            {6'd35, 6'd14}: alive_out = 1;
            {6'd35, 6'd15}: alive_out = 1;
            {6'd35, 6'd16}: alive_out = 1;
            {6'd35, 6'd17}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd35, 6'd20}: alive_out = 1;
            {6'd35, 6'd21}: alive_out = 1;
            {6'd35, 6'd22}: alive_out = 1;
            {6'd35, 6'd23}: alive_out = 1;
            {6'd35, 6'd24}: alive_out = 1;
            {6'd35, 6'd25}: alive_out = 1;
            {6'd35, 6'd26}: alive_out = 1;
            {6'd35, 6'd27}: alive_out = 1;
            {6'd35, 6'd28}: alive_out = 1;
            {6'd35, 6'd29}: alive_out = 1;
            {6'd35, 6'd30}: alive_out = 1;
            {6'd35, 6'd31}: alive_out = 1;
            {6'd35, 6'd32}: alive_out = 1;
            {6'd35, 6'd33}: alive_out = 1;
            {6'd35, 6'd34}: alive_out = 1;
            {6'd35, 6'd35}: alive_out = 1;
            {6'd35, 6'd36}: alive_out = 1;
            {6'd35, 6'd37}: alive_out = 1;
            {6'd35, 6'd38}: alive_out = 1;
            {6'd35, 6'd39}: alive_out = 1;
            {6'd35, 6'd40}: alive_out = 1;
            {6'd35, 6'd41}: alive_out = 1;
            {6'd35, 6'd42}: alive_out = 1;
            {6'd35, 6'd43}: alive_out = 1;
            {6'd35, 6'd44}: alive_out = 1;
            {6'd35, 6'd45}: alive_out = 1;
            {6'd35, 6'd46}: alive_out = 1;
            {6'd38, 6'd2}: alive_out = 1;
            {6'd38, 6'd3}: alive_out = 1;
            {6'd38, 6'd4}: alive_out = 1;
            {6'd38, 6'd5}: alive_out = 1;
            {6'd38, 6'd6}: alive_out = 1;
            {6'd38, 6'd7}: alive_out = 1;
            {6'd38, 6'd8}: alive_out = 1;
            {6'd38, 6'd9}: alive_out = 1;
            {6'd38, 6'd10}: alive_out = 1;
            {6'd38, 6'd11}: alive_out = 1;
            {6'd38, 6'd12}: alive_out = 1;
            {6'd38, 6'd13}: alive_out = 1;
            {6'd38, 6'd14}: alive_out = 1;
            {6'd38, 6'd15}: alive_out = 1;
            {6'd38, 6'd16}: alive_out = 1;
            {6'd38, 6'd17}: alive_out = 1;
            {6'd38, 6'd18}: alive_out = 1;
            {6'd38, 6'd19}: alive_out = 1;
            {6'd38, 6'd20}: alive_out = 1;
            {6'd38, 6'd21}: alive_out = 1;
            {6'd38, 6'd22}: alive_out = 1;
            {6'd38, 6'd23}: alive_out = 1;
            {6'd38, 6'd24}: alive_out = 1;
            {6'd38, 6'd25}: alive_out = 1;
            {6'd38, 6'd26}: alive_out = 1;
            {6'd38, 6'd27}: alive_out = 1;
            {6'd38, 6'd28}: alive_out = 1;
            {6'd38, 6'd29}: alive_out = 1;
            {6'd38, 6'd30}: alive_out = 1;
            {6'd38, 6'd31}: alive_out = 1;
            {6'd38, 6'd32}: alive_out = 1;
            {6'd38, 6'd33}: alive_out = 1;
            {6'd38, 6'd34}: alive_out = 1;
            {6'd38, 6'd35}: alive_out = 1;
            {6'd38, 6'd36}: alive_out = 1;
            {6'd38, 6'd37}: alive_out = 1;
            {6'd38, 6'd38}: alive_out = 1;
            {6'd38, 6'd39}: alive_out = 1;
            {6'd38, 6'd40}: alive_out = 1;
            {6'd38, 6'd41}: alive_out = 1;
            {6'd38, 6'd42}: alive_out = 1;
            {6'd38, 6'd43}: alive_out = 1;
            {6'd38, 6'd44}: alive_out = 1;
            {6'd38, 6'd45}: alive_out = 1;
            {6'd38, 6'd46}: alive_out = 1;
            {6'd39, 6'd2}: alive_out = 1;
            {6'd39, 6'd3}: alive_out = 1;
            {6'd39, 6'd4}: alive_out = 1;
            {6'd39, 6'd5}: alive_out = 1;
            {6'd39, 6'd6}: alive_out = 1;
            {6'd39, 6'd7}: alive_out = 1;
            {6'd39, 6'd8}: alive_out = 1;
            {6'd39, 6'd9}: alive_out = 1;
            {6'd39, 6'd10}: alive_out = 1;
            {6'd39, 6'd11}: alive_out = 1;
            {6'd39, 6'd12}: alive_out = 1;
            {6'd39, 6'd13}: alive_out = 1;
            {6'd39, 6'd14}: alive_out = 1;
            {6'd39, 6'd15}: alive_out = 1;
            {6'd39, 6'd16}: alive_out = 1;
            {6'd39, 6'd17}: alive_out = 1;
            {6'd39, 6'd18}: alive_out = 1;
            {6'd39, 6'd19}: alive_out = 1;
            {6'd39, 6'd20}: alive_out = 1;
            {6'd39, 6'd21}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd39, 6'd23}: alive_out = 1;
            {6'd39, 6'd24}: alive_out = 1;
            {6'd39, 6'd25}: alive_out = 1;
            {6'd39, 6'd26}: alive_out = 1;
            {6'd39, 6'd27}: alive_out = 1;
            {6'd39, 6'd28}: alive_out = 1;
            {6'd39, 6'd29}: alive_out = 1;
            {6'd39, 6'd30}: alive_out = 1;
            {6'd39, 6'd31}: alive_out = 1;
            {6'd39, 6'd32}: alive_out = 1;
            {6'd39, 6'd33}: alive_out = 1;
            {6'd39, 6'd34}: alive_out = 1;
            {6'd39, 6'd35}: alive_out = 1;
            {6'd39, 6'd36}: alive_out = 1;
            {6'd39, 6'd37}: alive_out = 1;
            {6'd39, 6'd38}: alive_out = 1;
            {6'd39, 6'd39}: alive_out = 1;
            {6'd39, 6'd40}: alive_out = 1;
            {6'd39, 6'd41}: alive_out = 1;
            {6'd39, 6'd42}: alive_out = 1;
            {6'd39, 6'd43}: alive_out = 1;
            {6'd39, 6'd44}: alive_out = 1;
            {6'd39, 6'd45}: alive_out = 1;
            {6'd39, 6'd46}: alive_out = 1;
            {6'd42, 6'd2}: alive_out = 1;
            {6'd42, 6'd3}: alive_out = 1;
            {6'd42, 6'd4}: alive_out = 1;
            {6'd42, 6'd5}: alive_out = 1;
            {6'd42, 6'd6}: alive_out = 1;
            {6'd42, 6'd7}: alive_out = 1;
            {6'd42, 6'd8}: alive_out = 1;
            {6'd42, 6'd9}: alive_out = 1;
            {6'd42, 6'd10}: alive_out = 1;
            {6'd42, 6'd11}: alive_out = 1;
            {6'd42, 6'd12}: alive_out = 1;
            {6'd42, 6'd13}: alive_out = 1;
            {6'd42, 6'd14}: alive_out = 1;
            {6'd42, 6'd15}: alive_out = 1;
            {6'd42, 6'd16}: alive_out = 1;
            {6'd42, 6'd17}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd42, 6'd19}: alive_out = 1;
            {6'd42, 6'd20}: alive_out = 1;
            {6'd42, 6'd21}: alive_out = 1;
            {6'd42, 6'd22}: alive_out = 1;
            {6'd42, 6'd23}: alive_out = 1;
            {6'd42, 6'd24}: alive_out = 1;
            {6'd42, 6'd25}: alive_out = 1;
            {6'd42, 6'd26}: alive_out = 1;
            {6'd42, 6'd27}: alive_out = 1;
            {6'd42, 6'd28}: alive_out = 1;
            {6'd42, 6'd29}: alive_out = 1;
            {6'd42, 6'd30}: alive_out = 1;
            {6'd42, 6'd31}: alive_out = 1;
            {6'd42, 6'd32}: alive_out = 1;
            {6'd42, 6'd33}: alive_out = 1;
            {6'd42, 6'd34}: alive_out = 1;
            {6'd42, 6'd35}: alive_out = 1;
            {6'd42, 6'd36}: alive_out = 1;
            {6'd42, 6'd37}: alive_out = 1;
            {6'd42, 6'd38}: alive_out = 1;
            {6'd42, 6'd39}: alive_out = 1;
            {6'd42, 6'd40}: alive_out = 1;
            {6'd42, 6'd41}: alive_out = 1;
            {6'd42, 6'd42}: alive_out = 1;
            {6'd42, 6'd43}: alive_out = 1;
            {6'd42, 6'd44}: alive_out = 1;
            {6'd42, 6'd45}: alive_out = 1;
            {6'd42, 6'd46}: alive_out = 1;
            {6'd43, 6'd2}: alive_out = 1;
            {6'd43, 6'd3}: alive_out = 1;
            {6'd43, 6'd4}: alive_out = 1;
            {6'd43, 6'd5}: alive_out = 1;
            {6'd43, 6'd6}: alive_out = 1;
            {6'd43, 6'd7}: alive_out = 1;
            {6'd43, 6'd8}: alive_out = 1;
            {6'd43, 6'd9}: alive_out = 1;
            {6'd43, 6'd10}: alive_out = 1;
            {6'd43, 6'd11}: alive_out = 1;
            {6'd43, 6'd12}: alive_out = 1;
            {6'd43, 6'd13}: alive_out = 1;
            {6'd43, 6'd14}: alive_out = 1;
            {6'd43, 6'd15}: alive_out = 1;
            {6'd43, 6'd16}: alive_out = 1;
            {6'd43, 6'd17}: alive_out = 1;
            {6'd43, 6'd18}: alive_out = 1;
            {6'd43, 6'd19}: alive_out = 1;
            {6'd43, 6'd20}: alive_out = 1;
            {6'd43, 6'd21}: alive_out = 1;
            {6'd43, 6'd22}: alive_out = 1;
            {6'd43, 6'd23}: alive_out = 1;
            {6'd43, 6'd24}: alive_out = 1;
            {6'd43, 6'd25}: alive_out = 1;
            {6'd43, 6'd26}: alive_out = 1;
            {6'd43, 6'd27}: alive_out = 1;
            {6'd43, 6'd28}: alive_out = 1;
            {6'd43, 6'd29}: alive_out = 1;
            {6'd43, 6'd30}: alive_out = 1;
            {6'd43, 6'd31}: alive_out = 1;
            {6'd43, 6'd32}: alive_out = 1;
            {6'd43, 6'd33}: alive_out = 1;
            {6'd43, 6'd34}: alive_out = 1;
            {6'd43, 6'd35}: alive_out = 1;
            {6'd43, 6'd36}: alive_out = 1;
            {6'd43, 6'd37}: alive_out = 1;
            {6'd43, 6'd38}: alive_out = 1;
            {6'd43, 6'd39}: alive_out = 1;
            {6'd43, 6'd40}: alive_out = 1;
            {6'd43, 6'd41}: alive_out = 1;
            {6'd43, 6'd42}: alive_out = 1;
            {6'd43, 6'd43}: alive_out = 1;
            {6'd43, 6'd44}: alive_out = 1;
            {6'd43, 6'd45}: alive_out = 1;
            {6'd43, 6'd46}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module trafficcircle(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd1, 6'd20}: alive_out = 1;
            {6'd1, 6'd21}: alive_out = 1;
            {6'd1, 6'd26}: alive_out = 1;
            {6'd1, 6'd27}: alive_out = 1;
            {6'd2, 6'd20}: alive_out = 1;
            {6'd2, 6'd22}: alive_out = 1;
            {6'd2, 6'd25}: alive_out = 1;
            {6'd2, 6'd27}: alive_out = 1;
            {6'd3, 6'd22}: alive_out = 1;
            {6'd3, 6'd25}: alive_out = 1;
            {6'd4, 6'd21}: alive_out = 1;
            {6'd4, 6'd22}: alive_out = 1;
            {6'd4, 6'd25}: alive_out = 1;
            {6'd4, 6'd26}: alive_out = 1;
            {6'd5, 6'd20}: alive_out = 1;
            {6'd5, 6'd21}: alive_out = 1;
            {6'd5, 6'd22}: alive_out = 1;
            {6'd5, 6'd25}: alive_out = 1;
            {6'd5, 6'd26}: alive_out = 1;
            {6'd5, 6'd27}: alive_out = 1;
            {6'd6, 6'd22}: alive_out = 1;
            {6'd6, 6'd25}: alive_out = 1;
            {6'd7, 6'd16}: alive_out = 1;
            {6'd7, 6'd17}: alive_out = 1;
            {6'd8, 6'd15}: alive_out = 1;
            {6'd8, 6'd16}: alive_out = 1;
            {6'd8, 6'd17}: alive_out = 1;
            {6'd9, 6'd14}: alive_out = 1;
            {6'd9, 6'd16}: alive_out = 1;
            {6'd9, 6'd17}: alive_out = 1;
            {6'd10, 6'd13}: alive_out = 1;
            {6'd10, 6'd15}: alive_out = 1;
            {6'd11, 6'd13}: alive_out = 1;
            {6'd11, 6'd16}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd11, 6'd22}: alive_out = 1;
            {6'd11, 6'd23}: alive_out = 1;
            {6'd12, 6'd14}: alive_out = 1;
            {6'd12, 6'd15}: alive_out = 1;
            {6'd13, 6'd19}: alive_out = 1;
            {6'd13, 6'd25}: alive_out = 1;
            {6'd13, 6'd38}: alive_out = 1;
            {6'd13, 6'd39}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd25}: alive_out = 1;
            {6'd14, 6'd37}: alive_out = 1;
            {6'd14, 6'd40}: alive_out = 1;
            {6'd15, 6'd19}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd15, 6'd37}: alive_out = 1;
            {6'd15, 6'd39}: alive_out = 1;
            {6'd15, 6'd42}: alive_out = 1;
            {6'd16, 6'd38}: alive_out = 1;
            {6'd17, 6'd21}: alive_out = 1;
            {6'd17, 6'd22}: alive_out = 1;
            {6'd17, 6'd23}: alive_out = 1;
            {6'd17, 6'd39}: alive_out = 1;
            {6'd17, 6'd40}: alive_out = 1;
            {6'd17, 6'd42}: alive_out = 1;
            {6'd18, 6'd41}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd20, 6'd24}: alive_out = 1;
            {6'd20, 6'd37}: alive_out = 1;
            {6'd20, 6'd44}: alive_out = 1;
            {6'd20, 6'd47}: alive_out = 1;
            {6'd20, 6'd48}: alive_out = 1;
            {6'd21, 6'd35}: alive_out = 1;
            {6'd21, 6'd44}: alive_out = 1;
            {6'd21, 6'd45}: alive_out = 1;
            {6'd21, 6'd48}: alive_out = 1;
            {6'd22, 6'd1}: alive_out = 1;
            {6'd22, 6'd2}: alive_out = 1;
            {6'd22, 6'd5}: alive_out = 1;
            {6'd22, 6'd20}: alive_out = 1;
            {6'd22, 6'd26}: alive_out = 1;
            {6'd22, 6'd35}: alive_out = 1;
            {6'd22, 6'd43}: alive_out = 1;
            {6'd22, 6'd44}: alive_out = 1;
            {6'd22, 6'd45}: alive_out = 1;
            {6'd22, 6'd46}: alive_out = 1;
            {6'd22, 6'd47}: alive_out = 1;
            {6'd23, 6'd1}: alive_out = 1;
            {6'd23, 6'd4}: alive_out = 1;
            {6'd23, 6'd5}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd23, 6'd37}: alive_out = 1;
            {6'd24, 6'd2}: alive_out = 1;
            {6'd24, 6'd3}: alive_out = 1;
            {6'd24, 6'd4}: alive_out = 1;
            {6'd24, 6'd5}: alive_out = 1;
            {6'd24, 6'd6}: alive_out = 1;
            {6'd24, 6'd14}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd26}: alive_out = 1;
            {6'd25, 6'd14}: alive_out = 1;
            {6'd25, 6'd43}: alive_out = 1;
            {6'd25, 6'd44}: alive_out = 1;
            {6'd25, 6'd45}: alive_out = 1;
            {6'd25, 6'd46}: alive_out = 1;
            {6'd25, 6'd47}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd44}: alive_out = 1;
            {6'd26, 6'd45}: alive_out = 1;
            {6'd26, 6'd48}: alive_out = 1;
            {6'd27, 6'd2}: alive_out = 1;
            {6'd27, 6'd3}: alive_out = 1;
            {6'd27, 6'd4}: alive_out = 1;
            {6'd27, 6'd5}: alive_out = 1;
            {6'd27, 6'd6}: alive_out = 1;
            {6'd27, 6'd10}: alive_out = 1;
            {6'd27, 6'd11}: alive_out = 1;
            {6'd27, 6'd12}: alive_out = 1;
            {6'd27, 6'd16}: alive_out = 1;
            {6'd27, 6'd17}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd44}: alive_out = 1;
            {6'd27, 6'd47}: alive_out = 1;
            {6'd27, 6'd48}: alive_out = 1;
            {6'd28, 6'd1}: alive_out = 1;
            {6'd28, 6'd4}: alive_out = 1;
            {6'd28, 6'd5}: alive_out = 1;
            {6'd29, 6'd1}: alive_out = 1;
            {6'd29, 6'd2}: alive_out = 1;
            {6'd29, 6'd5}: alive_out = 1;
            {6'd29, 6'd14}: alive_out = 1;
            {6'd30, 6'd14}: alive_out = 1;
            {6'd31, 6'd8}: alive_out = 1;
            {6'd31, 6'd10}: alive_out = 1;
            {6'd31, 6'd14}: alive_out = 1;
            {6'd32, 6'd7}: alive_out = 1;
            {6'd32, 6'd26}: alive_out = 1;
            {6'd32, 6'd27}: alive_out = 1;
            {6'd32, 6'd28}: alive_out = 1;
            {6'd33, 6'd8}: alive_out = 1;
            {6'd33, 6'd11}: alive_out = 1;
            {6'd34, 6'd8}: alive_out = 1;
            {6'd34, 6'd10}: alive_out = 1;
            {6'd34, 6'd12}: alive_out = 1;
            {6'd34, 6'd24}: alive_out = 1;
            {6'd34, 6'd30}: alive_out = 1;
            {6'd35, 6'd9}: alive_out = 1;
            {6'd35, 6'd12}: alive_out = 1;
            {6'd35, 6'd24}: alive_out = 1;
            {6'd35, 6'd30}: alive_out = 1;
            {6'd36, 6'd10}: alive_out = 1;
            {6'd36, 6'd11}: alive_out = 1;
            {6'd36, 6'd24}: alive_out = 1;
            {6'd36, 6'd30}: alive_out = 1;
            {6'd37, 6'd34}: alive_out = 1;
            {6'd37, 6'd35}: alive_out = 1;
            {6'd38, 6'd26}: alive_out = 1;
            {6'd38, 6'd27}: alive_out = 1;
            {6'd38, 6'd28}: alive_out = 1;
            {6'd38, 6'd33}: alive_out = 1;
            {6'd38, 6'd36}: alive_out = 1;
            {6'd39, 6'd32}: alive_out = 1;
            {6'd39, 6'd34}: alive_out = 1;
            {6'd39, 6'd36}: alive_out = 1;
            {6'd40, 6'd31}: alive_out = 1;
            {6'd40, 6'd32}: alive_out = 1;
            {6'd40, 6'd33}: alive_out = 1;
            {6'd40, 6'd35}: alive_out = 1;
            {6'd41, 6'd31}: alive_out = 1;
            {6'd41, 6'd32}: alive_out = 1;
            {6'd41, 6'd33}: alive_out = 1;
            {6'd43, 6'd24}: alive_out = 1;
            {6'd43, 6'd27}: alive_out = 1;
            {6'd44, 6'd22}: alive_out = 1;
            {6'd44, 6'd23}: alive_out = 1;
            {6'd44, 6'd24}: alive_out = 1;
            {6'd44, 6'd27}: alive_out = 1;
            {6'd44, 6'd28}: alive_out = 1;
            {6'd44, 6'd29}: alive_out = 1;
            {6'd45, 6'd23}: alive_out = 1;
            {6'd45, 6'd24}: alive_out = 1;
            {6'd45, 6'd27}: alive_out = 1;
            {6'd45, 6'd28}: alive_out = 1;
            {6'd46, 6'd24}: alive_out = 1;
            {6'd46, 6'd27}: alive_out = 1;
            {6'd47, 6'd22}: alive_out = 1;
            {6'd47, 6'd24}: alive_out = 1;
            {6'd47, 6'd27}: alive_out = 1;
            {6'd47, 6'd29}: alive_out = 1;
            {6'd48, 6'd22}: alive_out = 1;
            {6'd48, 6'd23}: alive_out = 1;
            {6'd48, 6'd28}: alive_out = 1;
            {6'd48, 6'd29}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module superfountain(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd2, 6'd24}: alive_out = 1;
            {6'd5, 6'd15}: alive_out = 1;
            {6'd5, 6'd21}: alive_out = 1;
            {6'd5, 6'd27}: alive_out = 1;
            {6'd5, 6'd33}: alive_out = 1;
            {6'd6, 6'd14}: alive_out = 1;
            {6'd6, 6'd16}: alive_out = 1;
            {6'd6, 6'd17}: alive_out = 1;
            {6'd6, 6'd18}: alive_out = 1;
            {6'd6, 6'd20}: alive_out = 1;
            {6'd6, 6'd22}: alive_out = 1;
            {6'd6, 6'd23}: alive_out = 1;
            {6'd6, 6'd24}: alive_out = 1;
            {6'd6, 6'd25}: alive_out = 1;
            {6'd6, 6'd26}: alive_out = 1;
            {6'd6, 6'd28}: alive_out = 1;
            {6'd6, 6'd30}: alive_out = 1;
            {6'd6, 6'd31}: alive_out = 1;
            {6'd6, 6'd32}: alive_out = 1;
            {6'd6, 6'd34}: alive_out = 1;
            {6'd7, 6'd15}: alive_out = 1;
            {6'd7, 6'd18}: alive_out = 1;
            {6'd7, 6'd23}: alive_out = 1;
            {6'd7, 6'd25}: alive_out = 1;
            {6'd7, 6'd30}: alive_out = 1;
            {6'd7, 6'd33}: alive_out = 1;
            {6'd8, 6'd18}: alive_out = 1;
            {6'd8, 6'd23}: alive_out = 1;
            {6'd8, 6'd25}: alive_out = 1;
            {6'd8, 6'd30}: alive_out = 1;
            {6'd10, 6'd19}: alive_out = 1;
            {6'd10, 6'd20}: alive_out = 1;
            {6'd10, 6'd22}: alive_out = 1;
            {6'd10, 6'd23}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd10, 6'd26}: alive_out = 1;
            {6'd10, 6'd28}: alive_out = 1;
            {6'd10, 6'd29}: alive_out = 1;
            {6'd11, 6'd13}: alive_out = 1;
            {6'd11, 6'd14}: alive_out = 1;
            {6'd11, 6'd19}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd11, 6'd22}: alive_out = 1;
            {6'd11, 6'd23}: alive_out = 1;
            {6'd11, 6'd25}: alive_out = 1;
            {6'd11, 6'd26}: alive_out = 1;
            {6'd11, 6'd27}: alive_out = 1;
            {6'd11, 6'd29}: alive_out = 1;
            {6'd11, 6'd34}: alive_out = 1;
            {6'd11, 6'd35}: alive_out = 1;
            {6'd12, 6'd13}: alive_out = 1;
            {6'd12, 6'd16}: alive_out = 1;
            {6'd12, 6'd18}: alive_out = 1;
            {6'd12, 6'd22}: alive_out = 1;
            {6'd12, 6'd26}: alive_out = 1;
            {6'd12, 6'd30}: alive_out = 1;
            {6'd12, 6'd32}: alive_out = 1;
            {6'd12, 6'd35}: alive_out = 1;
            {6'd13, 6'd14}: alive_out = 1;
            {6'd13, 6'd15}: alive_out = 1;
            {6'd13, 6'd21}: alive_out = 1;
            {6'd13, 6'd27}: alive_out = 1;
            {6'd13, 6'd33}: alive_out = 1;
            {6'd13, 6'd34}: alive_out = 1;
            {6'd14, 6'd17}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd23}: alive_out = 1;
            {6'd14, 6'd25}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd14, 6'd31}: alive_out = 1;
            {6'd15, 6'd14}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd15, 6'd16}: alive_out = 1;
            {6'd15, 6'd17}: alive_out = 1;
            {6'd15, 6'd23}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd15, 6'd31}: alive_out = 1;
            {6'd15, 6'd32}: alive_out = 1;
            {6'd15, 6'd33}: alive_out = 1;
            {6'd15, 6'd34}: alive_out = 1;
            {6'd16, 6'd14}: alive_out = 1;
            {6'd16, 6'd17}: alive_out = 1;
            {6'd16, 6'd19}: alive_out = 1;
            {6'd16, 6'd24}: alive_out = 1;
            {6'd16, 6'd29}: alive_out = 1;
            {6'd16, 6'd31}: alive_out = 1;
            {6'd16, 6'd34}: alive_out = 1;
            {6'd17, 6'd12}: alive_out = 1;
            {6'd17, 6'd14}: alive_out = 1;
            {6'd17, 6'd17}: alive_out = 1;
            {6'd17, 6'd19}: alive_out = 1;
            {6'd17, 6'd20}: alive_out = 1;
            {6'd17, 6'd28}: alive_out = 1;
            {6'd17, 6'd29}: alive_out = 1;
            {6'd17, 6'd31}: alive_out = 1;
            {6'd17, 6'd34}: alive_out = 1;
            {6'd17, 6'd36}: alive_out = 1;
            {6'd18, 6'd12}: alive_out = 1;
            {6'd18, 6'd13}: alive_out = 1;
            {6'd18, 6'd18}: alive_out = 1;
            {6'd18, 6'd22}: alive_out = 1;
            {6'd18, 6'd23}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd18, 6'd26}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd18, 6'd35}: alive_out = 1;
            {6'd18, 6'd36}: alive_out = 1;
            {6'd19, 6'd19}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd19, 6'd21}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd19, 6'd28}: alive_out = 1;
            {6'd19, 6'd29}: alive_out = 1;
            {6'd20, 6'd16}: alive_out = 1;
            {6'd20, 6'd17}: alive_out = 1;
            {6'd20, 6'd18}: alive_out = 1;
            {6'd20, 6'd24}: alive_out = 1;
            {6'd21, 6'd15}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd23}: alive_out = 1;
            {6'd21, 6'd24}: alive_out = 1;
            {6'd21, 6'd25}: alive_out = 1;
            {6'd21, 6'd29}: alive_out = 1;
            {6'd21, 6'd30}: alive_out = 1;
            {6'd21, 6'd31}: alive_out = 1;
            {6'd22, 6'd14}: alive_out = 1;
            {6'd22, 6'd16}: alive_out = 1;
            {6'd22, 6'd17}: alive_out = 1;
            {6'd22, 6'd19}: alive_out = 1;
            {6'd22, 6'd23}: alive_out = 1;
            {6'd22, 6'd26}: alive_out = 1;
            {6'd22, 6'd28}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd17}: alive_out = 1;
            {6'd23, 6'd18}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd21}: alive_out = 1;
            {6'd23, 6'd22}: alive_out = 1;
            {6'd23, 6'd23}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd30}: alive_out = 1;
            {6'd23, 6'd31}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd24, 6'd15}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd23}: alive_out = 1;
            {6'd24, 6'd24}: alive_out = 1;
            {6'd24, 6'd28}: alive_out = 1;
            {6'd24, 6'd31}: alive_out = 1;
            {6'd24, 6'd33}: alive_out = 1;
            {6'd24, 6'd34}: alive_out = 1;
            {6'd25, 6'd12}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd25, 6'd14}: alive_out = 1;
            {6'd25, 6'd21}: alive_out = 1;
            {6'd25, 6'd25}: alive_out = 1;
            {6'd25, 6'd27}: alive_out = 1;
            {6'd25, 6'd29}: alive_out = 1;
            {6'd25, 6'd31}: alive_out = 1;
            {6'd26, 6'd12}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd26}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd26, 6'd31}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd20}: alive_out = 1;
            {6'd27, 6'd21}: alive_out = 1;
            {6'd27, 6'd23}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd27, 6'd32}: alive_out = 1;
            {6'd27, 6'd33}: alive_out = 1;
            {6'd28, 6'd17}: alive_out = 1;
            {6'd28, 6'd18}: alive_out = 1;
            {6'd28, 6'd19}: alive_out = 1;
            {6'd28, 6'd21}: alive_out = 1;
            {6'd28, 6'd28}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd28, 6'd33}: alive_out = 1;
            {6'd29, 6'd16}: alive_out = 1;
            {6'd29, 6'd18}: alive_out = 1;
            {6'd29, 6'd21}: alive_out = 1;
            {6'd29, 6'd23}: alive_out = 1;
            {6'd29, 6'd24}: alive_out = 1;
            {6'd29, 6'd27}: alive_out = 1;
            {6'd29, 6'd28}: alive_out = 1;
            {6'd29, 6'd30}: alive_out = 1;
            {6'd29, 6'd31}: alive_out = 1;
            {6'd30, 6'd16}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd31, 6'd13}: alive_out = 1;
            {6'd31, 6'd14}: alive_out = 1;
            {6'd31, 6'd16}: alive_out = 1;
            {6'd31, 6'd19}: alive_out = 1;
            {6'd31, 6'd20}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd16}: alive_out = 1;
            {6'd32, 6'd18}: alive_out = 1;
            {6'd32, 6'd20}: alive_out = 1;
            {6'd32, 6'd23}: alive_out = 1;
            {6'd33, 6'd12}: alive_out = 1;
            {6'd33, 6'd15}: alive_out = 1;
            {6'd33, 6'd17}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd34, 6'd12}: alive_out = 1;
            {6'd34, 6'd13}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd34, 6'd22}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd34, 6'd25}: alive_out = 1;
            {6'd35, 6'd15}: alive_out = 1;
            {6'd35, 6'd16}: alive_out = 1;
            {6'd35, 6'd17}: alive_out = 1;
            {6'd35, 6'd22}: alive_out = 1;
            {6'd35, 6'd25}: alive_out = 1;
            {6'd36, 6'd15}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd36, 6'd19}: alive_out = 1;
            {6'd36, 6'd22}: alive_out = 1;
            {6'd36, 6'd23}: alive_out = 1;
            {6'd36, 6'd24}: alive_out = 1;
            {6'd37, 6'd12}: alive_out = 1;
            {6'd37, 6'd13}: alive_out = 1;
            {6'd37, 6'd15}: alive_out = 1;
            {6'd37, 6'd17}: alive_out = 1;
            {6'd38, 6'd12}: alive_out = 1;
            {6'd38, 6'd14}: alive_out = 1;
            {6'd39, 6'd14}: alive_out = 1;
            {6'd39, 6'd16}: alive_out = 1;
            {6'd39, 6'd18}: alive_out = 1;
            {6'd39, 6'd20}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd39, 6'd23}: alive_out = 1;
            {6'd39, 6'd24}: alive_out = 1;
            {6'd40, 6'd13}: alive_out = 1;
            {6'd40, 6'd14}: alive_out = 1;
            {6'd40, 6'd16}: alive_out = 1;
            {6'd40, 6'd18}: alive_out = 1;
            {6'd40, 6'd20}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;
            {6'd40, 6'd25}: alive_out = 1;
            {6'd41, 6'd17}: alive_out = 1;
            {6'd41, 6'd23}: alive_out = 1;
            {6'd41, 6'd25}: alive_out = 1;
            {6'd42, 6'd13}: alive_out = 1;
            {6'd42, 6'd14}: alive_out = 1;
            {6'd42, 6'd15}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd42, 6'd20}: alive_out = 1;
            {6'd42, 6'd21}: alive_out = 1;
            {6'd42, 6'd23}: alive_out = 1;
            {6'd42, 6'd24}: alive_out = 1;
            {6'd43, 6'd13}: alive_out = 1;
            {6'd43, 6'd16}: alive_out = 1;
            {6'd43, 6'd17}: alive_out = 1;
            {6'd43, 6'd19}: alive_out = 1;
            {6'd43, 6'd21}: alive_out = 1;
            {6'd44, 6'd14}: alive_out = 1;
            {6'd44, 6'd18}: alive_out = 1;
            {6'd44, 6'd19}: alive_out = 1;
            {6'd44, 6'd21}: alive_out = 1;
            {6'd45, 6'd15}: alive_out = 1;
            {6'd45, 6'd16}: alive_out = 1;
            {6'd45, 6'd20}: alive_out = 1;
            {6'd46, 6'd17}: alive_out = 1;
            {6'd46, 6'd18}: alive_out = 1;
            {6'd46, 6'd19}: alive_out = 1;
            {6'd47, 6'd17}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module harvester(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd16, 6'd29}: alive_out = 1;
            {6'd16, 6'd30}: alive_out = 1;
            {6'd16, 6'd31}: alive_out = 1;
            {6'd17, 6'd29}: alive_out = 1;
            {6'd17, 6'd30}: alive_out = 1;
            {6'd18, 6'd29}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd18, 6'd31}: alive_out = 1;
            {6'd19, 6'd29}: alive_out = 1;
            {6'd19, 6'd30}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd20, 6'd29}: alive_out = 1;
            {6'd21, 6'd28}: alive_out = 1;
            {6'd22, 6'd27}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd24, 6'd25}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd28, 6'd21}: alive_out = 1;
            {6'd29, 6'd20}: alive_out = 1;
            {6'd30, 6'd19}: alive_out = 1;
            {6'd31, 6'd18}: alive_out = 1;
            {6'd32, 6'd17}: alive_out = 1;
            {6'd33, 6'd17}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module wickstrecher(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd0, 6'd22}: alive_out = 1;
            {6'd1, 6'd20}: alive_out = 1;
            {6'd1, 6'd21}: alive_out = 1;
            {6'd1, 6'd22}: alive_out = 1;
            {6'd1, 6'd23}: alive_out = 1;
            {6'd1, 6'd24}: alive_out = 1;
            {6'd2, 6'd19}: alive_out = 1;
            {6'd2, 6'd25}: alive_out = 1;
            {6'd3, 6'd20}: alive_out = 1;
            {6'd3, 6'd21}: alive_out = 1;
            {6'd3, 6'd22}: alive_out = 1;
            {6'd3, 6'd24}: alive_out = 1;
            {6'd3, 6'd26}: alive_out = 1;
            {6'd4, 6'd22}: alive_out = 1;
            {6'd4, 6'd24}: alive_out = 1;
            {6'd4, 6'd26}: alive_out = 1;
            {6'd5, 6'd27}: alive_out = 1;
            {6'd5, 6'd28}: alive_out = 1;
            {6'd6, 6'd20}: alive_out = 1;
            {6'd6, 6'd21}: alive_out = 1;
            {6'd6, 6'd22}: alive_out = 1;
            {6'd6, 6'd23}: alive_out = 1;
            {6'd6, 6'd25}: alive_out = 1;
            {6'd6, 6'd27}: alive_out = 1;
            {6'd7, 6'd19}: alive_out = 1;
            {6'd7, 6'd23}: alive_out = 1;
            {6'd7, 6'd24}: alive_out = 1;
            {6'd7, 6'd25}: alive_out = 1;
            {6'd7, 6'd28}: alive_out = 1;
            {6'd8, 6'd19}: alive_out = 1;
            {6'd8, 6'd21}: alive_out = 1;
            {6'd8, 6'd22}: alive_out = 1;
            {6'd8, 6'd25}: alive_out = 1;
            {6'd8, 6'd26}: alive_out = 1;
            {6'd8, 6'd27}: alive_out = 1;
            {6'd8, 6'd28}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd9, 6'd19}: alive_out = 1;
            {6'd9, 6'd21}: alive_out = 1;
            {6'd10, 6'd17}: alive_out = 1;
            {6'd10, 6'd22}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd10, 6'd26}: alive_out = 1;
            {6'd10, 6'd27}: alive_out = 1;
            {6'd10, 6'd28}: alive_out = 1;
            {6'd11, 6'd18}: alive_out = 1;
            {6'd11, 6'd19}: alive_out = 1;
            {6'd11, 6'd20}: alive_out = 1;
            {6'd11, 6'd22}: alive_out = 1;
            {6'd11, 6'd24}: alive_out = 1;
            {6'd11, 6'd27}: alive_out = 1;
            {6'd11, 6'd29}: alive_out = 1;
            {6'd12, 6'd20}: alive_out = 1;
            {6'd12, 6'd23}: alive_out = 1;
            {6'd12, 6'd25}: alive_out = 1;
            {6'd12, 6'd29}: alive_out = 1;
            {6'd13, 6'd21}: alive_out = 1;
            {6'd13, 6'd23}: alive_out = 1;
            {6'd13, 6'd24}: alive_out = 1;
            {6'd13, 6'd26}: alive_out = 1;
            {6'd13, 6'd27}: alive_out = 1;
            {6'd13, 6'd28}: alive_out = 1;
            {6'd15, 6'd24}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd15, 6'd27}: alive_out = 1;
            {6'd15, 6'd28}: alive_out = 1;
            {6'd16, 6'd20}: alive_out = 1;
            {6'd16, 6'd24}: alive_out = 1;
            {6'd16, 6'd28}: alive_out = 1;
            {6'd17, 6'd19}: alive_out = 1;
            {6'd17, 6'd21}: alive_out = 1;
            {6'd17, 6'd23}: alive_out = 1;
            {6'd18, 6'd20}: alive_out = 1;
            {6'd19, 6'd23}: alive_out = 1;
            {6'd19, 6'd24}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd20, 6'd25}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd29}: alive_out = 1;
            {6'd21, 6'd24}: alive_out = 1;
            {6'd21, 6'd28}: alive_out = 1;
            {6'd21, 6'd29}: alive_out = 1;
            {6'd22, 6'd24}: alive_out = 1;
            {6'd24, 6'd24}: alive_out = 1;
            {6'd24, 6'd25}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd25, 6'd25}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd21}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd28}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd27, 6'd21}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd28, 6'd20}: alive_out = 1;
            {6'd28, 6'd21}: alive_out = 1;
            {6'd28, 6'd28}: alive_out = 1;
            {6'd28, 6'd29}: alive_out = 1;
            {6'd29, 6'd18}: alive_out = 1;
            {6'd29, 6'd31}: alive_out = 1;
            {6'd30, 6'd17}: alive_out = 1;
            {6'd30, 6'd20}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd29}: alive_out = 1;
            {6'd30, 6'd32}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd20}: alive_out = 1;
            {6'd31, 6'd22}: alive_out = 1;
            {6'd31, 6'd24}: alive_out = 1;
            {6'd31, 6'd25}: alive_out = 1;
            {6'd31, 6'd27}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd31, 6'd32}: alive_out = 1;
            {6'd32, 6'd19}: alive_out = 1;
            {6'd32, 6'd20}: alive_out = 1;
            {6'd32, 6'd29}: alive_out = 1;
            {6'd32, 6'd30}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd33, 6'd24}: alive_out = 1;
            {6'd33, 6'd25}: alive_out = 1;
            {6'd33, 6'd29}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd19}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd34, 6'd26}: alive_out = 1;
            {6'd34, 6'd30}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd35, 6'd30}: alive_out = 1;
            {6'd35, 6'd31}: alive_out = 1;
            {6'd36, 6'd19}: alive_out = 1;
            {6'd36, 6'd22}: alive_out = 1;
            {6'd36, 6'd27}: alive_out = 1;
            {6'd36, 6'd30}: alive_out = 1;
            {6'd37, 6'd20}: alive_out = 1;
            {6'd37, 6'd22}: alive_out = 1;
            {6'd37, 6'd27}: alive_out = 1;
            {6'd37, 6'd29}: alive_out = 1;
            {6'd39, 6'd21}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd39, 6'd27}: alive_out = 1;
            {6'd39, 6'd28}: alive_out = 1;
            {6'd40, 6'd22}: alive_out = 1;
            {6'd40, 6'd27}: alive_out = 1;
            {6'd41, 6'd20}: alive_out = 1;
            {6'd41, 6'd29}: alive_out = 1;
            {6'd42, 6'd20}: alive_out = 1;
            {6'd42, 6'd21}: alive_out = 1;
            {6'd42, 6'd23}: alive_out = 1;
            {6'd42, 6'd26}: alive_out = 1;
            {6'd42, 6'd28}: alive_out = 1;
            {6'd42, 6'd29}: alive_out = 1;
            {6'd43, 6'd21}: alive_out = 1;
            {6'd43, 6'd24}: alive_out = 1;
            {6'd43, 6'd25}: alive_out = 1;
            {6'd43, 6'd28}: alive_out = 1;
            {6'd45, 6'd20}: alive_out = 1;
            {6'd45, 6'd22}: alive_out = 1;
            {6'd45, 6'd27}: alive_out = 1;
            {6'd45, 6'd29}: alive_out = 1;
            {6'd46, 6'd20}: alive_out = 1;
            {6'd46, 6'd22}: alive_out = 1;
            {6'd46, 6'd27}: alive_out = 1;
            {6'd46, 6'd29}: alive_out = 1;
            {6'd48, 6'd20}: alive_out = 1;
            {6'd48, 6'd21}: alive_out = 1;
            {6'd48, 6'd22}: alive_out = 1;
            {6'd48, 6'd27}: alive_out = 1;
            {6'd48, 6'd28}: alive_out = 1;
            {6'd48, 6'd29}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module rectifier(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd4, 6'd17}: alive_out = 1;
            {6'd5, 6'd8}: alive_out = 1;
            {6'd5, 6'd15}: alive_out = 1;
            {6'd5, 6'd16}: alive_out = 1;
            {6'd5, 6'd17}: alive_out = 1;
            {6'd6, 6'd9}: alive_out = 1;
            {6'd6, 6'd10}: alive_out = 1;
            {6'd6, 6'd14}: alive_out = 1;
            {6'd7, 6'd8}: alive_out = 1;
            {6'd7, 6'd9}: alive_out = 1;
            {6'd7, 6'd14}: alive_out = 1;
            {6'd7, 6'd15}: alive_out = 1;
            {6'd13, 6'd24}: alive_out = 1;
            {6'd14, 6'd9}: alive_out = 1;
            {6'd14, 6'd10}: alive_out = 1;
            {6'd14, 6'd22}: alive_out = 1;
            {6'd14, 6'd23}: alive_out = 1;
            {6'd14, 6'd24}: alive_out = 1;
            {6'd15, 6'd8}: alive_out = 1;
            {6'd15, 6'd11}: alive_out = 1;
            {6'd15, 6'd21}: alive_out = 1;
            {6'd16, 6'd9}: alive_out = 1;
            {6'd16, 6'd10}: alive_out = 1;
            {6'd16, 6'd21}: alive_out = 1;
            {6'd16, 6'd22}: alive_out = 1;
            {6'd24, 6'd12}: alive_out = 1;
            {6'd24, 6'd13}: alive_out = 1;
            {6'd25, 6'd12}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd34, 6'd19}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd21}: alive_out = 1;
            {6'd35, 6'd24}: alive_out = 1;
            {6'd35, 6'd25}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd36, 6'd25}: alive_out = 1;
            {6'd37, 6'd19}: alive_out = 1;
            {6'd37, 6'd25}: alive_out = 1;
            {6'd37, 6'd26}: alive_out = 1;
            {6'd37, 6'd27}: alive_out = 1;
            {6'd38, 6'd22}: alive_out = 1;
            {6'd38, 6'd23}: alive_out = 1;
            {6'd38, 6'd25}: alive_out = 1;
            {6'd38, 6'd26}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd39, 6'd25}: alive_out = 1;
            {6'd39, 6'd27}: alive_out = 1;
            {6'd40, 6'd19}: alive_out = 1;
            {6'd40, 6'd24}: alive_out = 1;
            {6'd40, 6'd26}: alive_out = 1;
            {6'd40, 6'd27}: alive_out = 1;
            {6'd41, 6'd19}: alive_out = 1;
            {6'd41, 6'd20}: alive_out = 1;
            {6'd41, 6'd21}: alive_out = 1;
            {6'd41, 6'd22}: alive_out = 1;
            {6'd41, 6'd23}: alive_out = 1;
            {6'd43, 6'd21}: alive_out = 1;
            {6'd43, 6'd22}: alive_out = 1;
            {6'd43, 6'd24}: alive_out = 1;
            {6'd44, 6'd21}: alive_out = 1;
            {6'd44, 6'd23}: alive_out = 1;
            {6'd44, 6'd24}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module fly(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd20}: alive_out = 1;
            {6'd9, 6'd16}: alive_out = 1;
            {6'd9, 6'd17}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd9, 6'd20}: alive_out = 1;
            {6'd9, 6'd21}: alive_out = 1;
            {6'd9, 6'd22}: alive_out = 1;
            {6'd10, 6'd15}: alive_out = 1;
            {6'd10, 6'd22}: alive_out = 1;
            {6'd10, 6'd23}: alive_out = 1;
            {6'd11, 6'd16}: alive_out = 1;
            {6'd11, 6'd17}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd11, 6'd24}: alive_out = 1;
            {6'd11, 6'd28}: alive_out = 1;
            {6'd12, 6'd26}: alive_out = 1;
            {6'd12, 6'd27}: alive_out = 1;
            {6'd12, 6'd28}: alive_out = 1;
            {6'd12, 6'd29}: alive_out = 1;
            {6'd13, 6'd26}: alive_out = 1;
            {6'd13, 6'd30}: alive_out = 1;
            {6'd14, 6'd24}: alive_out = 1;
            {6'd14, 6'd27}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd15, 6'd25}: alive_out = 1;
            {6'd17, 6'd25}: alive_out = 1;
            {6'd17, 6'd26}: alive_out = 1;
            {6'd18, 6'd23}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd18, 6'd26}: alive_out = 1;
            {6'd18, 6'd27}: alive_out = 1;
            {6'd18, 6'd28}: alive_out = 1;
            {6'd19, 6'd19}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd19, 6'd22}: alive_out = 1;
            {6'd19, 6'd29}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd20, 6'd19}: alive_out = 1;
            {6'd20, 6'd20}: alive_out = 1;
            {6'd20, 6'd31}: alive_out = 1;
            {6'd20, 6'd32}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd21}: alive_out = 1;
            {6'd21, 6'd30}: alive_out = 1;
            {6'd21, 6'd32}: alive_out = 1;
            {6'd22, 6'd21}: alive_out = 1;
            {6'd22, 6'd22}: alive_out = 1;
            {6'd22, 6'd29}: alive_out = 1;
            {6'd22, 6'd30}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd21}: alive_out = 1;
            {6'd23, 6'd23}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd25}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd23, 6'd27}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd30}: alive_out = 1;
            {6'd23, 6'd31}: alive_out = 1;
            {6'd24, 6'd21}: alive_out = 1;
            {6'd24, 6'd30}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd31}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd26}: alive_out = 1;
            {6'd26, 6'd27}: alive_out = 1;
            {6'd26, 6'd28}: alive_out = 1;
            {6'd26, 6'd29}: alive_out = 1;
            {6'd26, 6'd31}: alive_out = 1;
            {6'd27, 6'd21}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd23}: alive_out = 1;
            {6'd27, 6'd24}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd27, 6'd26}: alive_out = 1;
            {6'd27, 6'd27}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd27, 6'd29}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd28, 6'd22}: alive_out = 1;
            {6'd28, 6'd24}: alive_out = 1;
            {6'd28, 6'd25}: alive_out = 1;
            {6'd28, 6'd26}: alive_out = 1;
            {6'd28, 6'd27}: alive_out = 1;
            {6'd28, 6'd29}: alive_out = 1;
            {6'd29, 6'd21}: alive_out = 1;
            {6'd29, 6'd25}: alive_out = 1;
            {6'd29, 6'd26}: alive_out = 1;
            {6'd29, 6'd30}: alive_out = 1;
            {6'd30, 6'd19}: alive_out = 1;
            {6'd30, 6'd20}: alive_out = 1;
            {6'd30, 6'd23}: alive_out = 1;
            {6'd30, 6'd24}: alive_out = 1;
            {6'd30, 6'd27}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd31}: alive_out = 1;
            {6'd30, 6'd32}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd32, 6'd21}: alive_out = 1;
            {6'd32, 6'd24}: alive_out = 1;
            {6'd32, 6'd27}: alive_out = 1;
            {6'd32, 6'd30}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd30}: alive_out = 1;
            {6'd33, 6'd31}: alive_out = 1;
            {6'd33, 6'd33}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd34, 6'd22}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd34, 6'd28}: alive_out = 1;
            {6'd34, 6'd29}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd34, 6'd33}: alive_out = 1;
            {6'd34, 6'd34}: alive_out = 1;
            {6'd35, 6'd20}: alive_out = 1;
            {6'd35, 6'd22}: alive_out = 1;
            {6'd35, 6'd25}: alive_out = 1;
            {6'd35, 6'd26}: alive_out = 1;
            {6'd35, 6'd29}: alive_out = 1;
            {6'd35, 6'd31}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd36, 6'd22}: alive_out = 1;
            {6'd36, 6'd29}: alive_out = 1;
            {6'd36, 6'd31}: alive_out = 1;
            {6'd36, 6'd33}: alive_out = 1;
            {6'd36, 6'd34}: alive_out = 1;
            {6'd37, 6'd23}: alive_out = 1;
            {6'd37, 6'd24}: alive_out = 1;
            {6'd37, 6'd27}: alive_out = 1;
            {6'd37, 6'd28}: alive_out = 1;
            {6'd38, 6'd18}: alive_out = 1;
            {6'd38, 6'd21}: alive_out = 1;
            {6'd38, 6'd24}: alive_out = 1;
            {6'd38, 6'd27}: alive_out = 1;
            {6'd38, 6'd30}: alive_out = 1;
            {6'd38, 6'd33}: alive_out = 1;
            {6'd39, 6'd21}: alive_out = 1;
            {6'd39, 6'd30}: alive_out = 1;
            {6'd40, 6'd17}: alive_out = 1;
            {6'd40, 6'd19}: alive_out = 1;
            {6'd40, 6'd32}: alive_out = 1;
            {6'd40, 6'd34}: alive_out = 1;
            {6'd41, 6'd18}: alive_out = 1;
            {6'd41, 6'd33}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module spacefiller(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd0, 6'd14}: alive_out = 1;
            {6'd0, 6'd15}: alive_out = 1;
            {6'd0, 6'd16}: alive_out = 1;
            {6'd0, 6'd22}: alive_out = 1;
            {6'd0, 6'd23}: alive_out = 1;
            {6'd0, 6'd24}: alive_out = 1;
            {6'd1, 6'd14}: alive_out = 1;
            {6'd1, 6'd17}: alive_out = 1;
            {6'd1, 6'd21}: alive_out = 1;
            {6'd1, 6'd24}: alive_out = 1;
            {6'd2, 6'd14}: alive_out = 1;
            {6'd2, 6'd24}: alive_out = 1;
            {6'd3, 6'd14}: alive_out = 1;
            {6'd3, 6'd24}: alive_out = 1;
            {6'd4, 6'd15}: alive_out = 1;
            {6'd4, 6'd17}: alive_out = 1;
            {6'd4, 6'd21}: alive_out = 1;
            {6'd4, 6'd23}: alive_out = 1;
            {6'd6, 6'd18}: alive_out = 1;
            {6'd6, 6'd19}: alive_out = 1;
            {6'd6, 6'd20}: alive_out = 1;
            {6'd7, 6'd17}: alive_out = 1;
            {6'd7, 6'd21}: alive_out = 1;
            {6'd8, 6'd17}: alive_out = 1;
            {6'd8, 6'd21}: alive_out = 1;
            {6'd9, 6'd16}: alive_out = 1;
            {6'd9, 6'd22}: alive_out = 1;
            {6'd11, 6'd17}: alive_out = 1;
            {6'd11, 6'd21}: alive_out = 1;
            {6'd12, 6'd18}: alive_out = 1;
            {6'd12, 6'd19}: alive_out = 1;
            {6'd12, 6'd20}: alive_out = 1;
            {6'd13, 6'd22}: alive_out = 1;
            {6'd14, 6'd21}: alive_out = 1;
            {6'd14, 6'd22}: alive_out = 1;
            {6'd14, 6'd23}: alive_out = 1;
            {6'd15, 6'd21}: alive_out = 1;
            {6'd15, 6'd23}: alive_out = 1;
            {6'd15, 6'd24}: alive_out = 1;
            {6'd16, 6'd24}: alive_out = 1;
            {6'd16, 6'd25}: alive_out = 1;
            {6'd17, 6'd24}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd19, 6'd13}: alive_out = 1;
            {6'd19, 6'd22}: alive_out = 1;
            {6'd19, 6'd24}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd27}: alive_out = 1;
            {6'd20, 6'd12}: alive_out = 1;
            {6'd20, 6'd18}: alive_out = 1;
            {6'd20, 6'd21}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd24}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd28}: alive_out = 1;
            {6'd20, 6'd30}: alive_out = 1;
            {6'd20, 6'd35}: alive_out = 1;
            {6'd20, 6'd36}: alive_out = 1;
            {6'd21, 6'd12}: alive_out = 1;
            {6'd21, 6'd18}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd20}: alive_out = 1;
            {6'd21, 6'd22}: alive_out = 1;
            {6'd21, 6'd24}: alive_out = 1;
            {6'd21, 6'd26}: alive_out = 1;
            {6'd21, 6'd28}: alive_out = 1;
            {6'd21, 6'd30}: alive_out = 1;
            {6'd21, 6'd33}: alive_out = 1;
            {6'd21, 6'd34}: alive_out = 1;
            {6'd21, 6'd36}: alive_out = 1;
            {6'd21, 6'd37}: alive_out = 1;
            {6'd22, 6'd12}: alive_out = 1;
            {6'd22, 6'd13}: alive_out = 1;
            {6'd22, 6'd14}: alive_out = 1;
            {6'd22, 6'd15}: alive_out = 1;
            {6'd22, 6'd16}: alive_out = 1;
            {6'd22, 6'd18}: alive_out = 1;
            {6'd22, 6'd20}: alive_out = 1;
            {6'd22, 6'd22}: alive_out = 1;
            {6'd22, 6'd24}: alive_out = 1;
            {6'd22, 6'd26}: alive_out = 1;
            {6'd22, 6'd28}: alive_out = 1;
            {6'd22, 6'd30}: alive_out = 1;
            {6'd22, 6'd31}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd22, 6'd34}: alive_out = 1;
            {6'd22, 6'd35}: alive_out = 1;
            {6'd22, 6'd36}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd22}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd33}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd22}: alive_out = 1;
            {6'd24, 6'd24}: alive_out = 1;
            {6'd24, 6'd26}: alive_out = 1;
            {6'd24, 6'd28}: alive_out = 1;
            {6'd24, 6'd29}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd22}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd25, 6'd26}: alive_out = 1;
            {6'd25, 6'd28}: alive_out = 1;
            {6'd25, 6'd33}: alive_out = 1;
            {6'd25, 6'd34}: alive_out = 1;
            {6'd25, 6'd35}: alive_out = 1;
            {6'd26, 6'd12}: alive_out = 1;
            {6'd26, 6'd13}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd15}: alive_out = 1;
            {6'd26, 6'd16}: alive_out = 1;
            {6'd26, 6'd18}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd24}: alive_out = 1;
            {6'd26, 6'd26}: alive_out = 1;
            {6'd26, 6'd28}: alive_out = 1;
            {6'd26, 6'd30}: alive_out = 1;
            {6'd26, 6'd31}: alive_out = 1;
            {6'd26, 6'd33}: alive_out = 1;
            {6'd26, 6'd34}: alive_out = 1;
            {6'd26, 6'd35}: alive_out = 1;
            {6'd26, 6'd36}: alive_out = 1;
            {6'd27, 6'd12}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd20}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd24}: alive_out = 1;
            {6'd27, 6'd26}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd27, 6'd33}: alive_out = 1;
            {6'd27, 6'd34}: alive_out = 1;
            {6'd27, 6'd36}: alive_out = 1;
            {6'd27, 6'd37}: alive_out = 1;
            {6'd28, 6'd12}: alive_out = 1;
            {6'd28, 6'd18}: alive_out = 1;
            {6'd28, 6'd21}: alive_out = 1;
            {6'd28, 6'd22}: alive_out = 1;
            {6'd28, 6'd24}: alive_out = 1;
            {6'd28, 6'd26}: alive_out = 1;
            {6'd28, 6'd28}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd28, 6'd35}: alive_out = 1;
            {6'd28, 6'd36}: alive_out = 1;
            {6'd29, 6'd13}: alive_out = 1;
            {6'd29, 6'd22}: alive_out = 1;
            {6'd29, 6'd24}: alive_out = 1;
            {6'd29, 6'd26}: alive_out = 1;
            {6'd29, 6'd27}: alive_out = 1;
            {6'd30, 6'd24}: alive_out = 1;
            {6'd30, 6'd25}: alive_out = 1;
            {6'd31, 6'd24}: alive_out = 1;
            {6'd32, 6'd24}: alive_out = 1;
            {6'd32, 6'd25}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd23}: alive_out = 1;
            {6'd33, 6'd24}: alive_out = 1;
            {6'd34, 6'd21}: alive_out = 1;
            {6'd34, 6'd22}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd35, 6'd22}: alive_out = 1;
            {6'd36, 6'd18}: alive_out = 1;
            {6'd36, 6'd19}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd37, 6'd17}: alive_out = 1;
            {6'd37, 6'd21}: alive_out = 1;
            {6'd39, 6'd16}: alive_out = 1;
            {6'd39, 6'd22}: alive_out = 1;
            {6'd40, 6'd17}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;
            {6'd41, 6'd17}: alive_out = 1;
            {6'd41, 6'd21}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd42, 6'd19}: alive_out = 1;
            {6'd42, 6'd20}: alive_out = 1;
            {6'd44, 6'd15}: alive_out = 1;
            {6'd44, 6'd17}: alive_out = 1;
            {6'd44, 6'd21}: alive_out = 1;
            {6'd44, 6'd23}: alive_out = 1;
            {6'd45, 6'd14}: alive_out = 1;
            {6'd45, 6'd24}: alive_out = 1;
            {6'd46, 6'd14}: alive_out = 1;
            {6'd46, 6'd24}: alive_out = 1;
            {6'd47, 6'd14}: alive_out = 1;
            {6'd47, 6'd17}: alive_out = 1;
            {6'd47, 6'd21}: alive_out = 1;
            {6'd47, 6'd24}: alive_out = 1;
            {6'd48, 6'd14}: alive_out = 1;
            {6'd48, 6'd15}: alive_out = 1;
            {6'd48, 6'd16}: alive_out = 1;
            {6'd48, 6'd22}: alive_out = 1;
            {6'd48, 6'd23}: alive_out = 1;
            {6'd48, 6'd24}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module pulsar(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd18, 6'd19}: alive_out = 1;
            {6'd18, 6'd20}: alive_out = 1;
            {6'd18, 6'd21}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd25}: alive_out = 1;
            {6'd18, 6'd26}: alive_out = 1;
            {6'd20, 6'd18}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd20, 6'd27}: alive_out = 1;
            {6'd21, 6'd18}: alive_out = 1;
            {6'd21, 6'd22}: alive_out = 1;
            {6'd21, 6'd23}: alive_out = 1;
            {6'd21, 6'd27}: alive_out = 1;
            {6'd22, 6'd18}: alive_out = 1;
            {6'd22, 6'd22}: alive_out = 1;
            {6'd22, 6'd23}: alive_out = 1;
            {6'd22, 6'd27}: alive_out = 1;
            {6'd23, 6'd19}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd21}: alive_out = 1;
            {6'd23, 6'd24}: alive_out = 1;
            {6'd23, 6'd25}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd25, 6'd19}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd21}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd25, 6'd25}: alive_out = 1;
            {6'd25, 6'd26}: alive_out = 1;
            {6'd26, 6'd18}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd26, 6'd27}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd23}: alive_out = 1;
            {6'd27, 6'd27}: alive_out = 1;
            {6'd28, 6'd18}: alive_out = 1;
            {6'd28, 6'd22}: alive_out = 1;
            {6'd28, 6'd23}: alive_out = 1;
            {6'd28, 6'd27}: alive_out = 1;
            {6'd30, 6'd19}: alive_out = 1;
            {6'd30, 6'd20}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd30, 6'd24}: alive_out = 1;
            {6'd30, 6'd25}: alive_out = 1;
            {6'd30, 6'd26}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module 10cellinfinitegrowth(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd21, 6'd27}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd23, 6'd27}: alive_out = 1;
            {6'd25, 6'd23}: alive_out = 1;
            {6'd25, 6'd24}: alive_out = 1;
            {6'd25, 6'd25}: alive_out = 1;
            {6'd27, 6'd22}: alive_out = 1;
            {6'd27, 6'd23}: alive_out = 1;
            {6'd27, 6'd24}: alive_out = 1;
            {6'd28, 6'd23}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module vacuumgun(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd0, 6'd7}: alive_out = 1;
            {6'd0, 6'd8}: alive_out = 1;
            {6'd0, 6'd14}: alive_out = 1;
            {6'd0, 6'd15}: alive_out = 1;
            {6'd1, 6'd3}: alive_out = 1;
            {6'd1, 6'd4}: alive_out = 1;
            {6'd1, 6'd7}: alive_out = 1;
            {6'd1, 6'd8}: alive_out = 1;
            {6'd1, 6'd14}: alive_out = 1;
            {6'd1, 6'd15}: alive_out = 1;
            {6'd1, 6'd18}: alive_out = 1;
            {6'd1, 6'd19}: alive_out = 1;
            {6'd2, 6'd3}: alive_out = 1;
            {6'd2, 6'd4}: alive_out = 1;
            {6'd2, 6'd18}: alive_out = 1;
            {6'd2, 6'd19}: alive_out = 1;
            {6'd14, 6'd40}: alive_out = 1;
            {6'd15, 6'd6}: alive_out = 1;
            {6'd15, 6'd7}: alive_out = 1;
            {6'd15, 6'd8}: alive_out = 1;
            {6'd15, 6'd14}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd15, 6'd16}: alive_out = 1;
            {6'd15, 6'd38}: alive_out = 1;
            {6'd15, 6'd39}: alive_out = 1;
            {6'd15, 6'd40}: alive_out = 1;
            {6'd16, 6'd6}: alive_out = 1;
            {6'd16, 6'd9}: alive_out = 1;
            {6'd16, 6'd10}: alive_out = 1;
            {6'd16, 6'd12}: alive_out = 1;
            {6'd16, 6'd13}: alive_out = 1;
            {6'd16, 6'd16}: alive_out = 1;
            {6'd16, 6'd37}: alive_out = 1;
            {6'd17, 6'd7}: alive_out = 1;
            {6'd17, 6'd8}: alive_out = 1;
            {6'd17, 6'd9}: alive_out = 1;
            {6'd17, 6'd13}: alive_out = 1;
            {6'd17, 6'd14}: alive_out = 1;
            {6'd17, 6'd15}: alive_out = 1;
            {6'd17, 6'd37}: alive_out = 1;
            {6'd17, 6'd38}: alive_out = 1;
            {6'd18, 6'd8}: alive_out = 1;
            {6'd18, 6'd14}: alive_out = 1;
            {6'd21, 6'd32}: alive_out = 1;
            {6'd21, 6'd33}: alive_out = 1;
            {6'd21, 6'd34}: alive_out = 1;
            {6'd21, 6'd36}: alive_out = 1;
            {6'd22, 6'd31}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd22, 6'd36}: alive_out = 1;
            {6'd22, 6'd37}: alive_out = 1;
            {6'd23, 6'd32}: alive_out = 1;
            {6'd23, 6'd33}: alive_out = 1;
            {6'd24, 6'd5}: alive_out = 1;
            {6'd24, 6'd6}: alive_out = 1;
            {6'd24, 6'd31}: alive_out = 1;
            {6'd24, 6'd38}: alive_out = 1;
            {6'd25, 6'd6}: alive_out = 1;
            {6'd25, 6'd35}: alive_out = 1;
            {6'd26, 6'd3}: alive_out = 1;
            {6'd26, 6'd4}: alive_out = 1;
            {6'd26, 6'd5}: alive_out = 1;
            {6'd26, 6'd37}: alive_out = 1;
            {6'd27, 6'd3}: alive_out = 1;
            {6'd27, 6'd35}: alive_out = 1;
            {6'd27, 6'd36}: alive_out = 1;
            {6'd27, 6'd37}: alive_out = 1;
            {6'd31, 6'd15}: alive_out = 1;
            {6'd31, 6'd16}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd22}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd17}: alive_out = 1;
            {6'd32, 6'd21}: alive_out = 1;
            {6'd32, 6'd24}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd20}: alive_out = 1;
            {6'd36, 6'd14}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd21}: alive_out = 1;
            {6'd36, 6'd24}: alive_out = 1;
            {6'd37, 6'd15}: alive_out = 1;
            {6'd37, 6'd23}: alive_out = 1;
            {6'd37, 6'd27}: alive_out = 1;
            {6'd37, 6'd28}: alive_out = 1;
            {6'd37, 6'd30}: alive_out = 1;
            {6'd37, 6'd34}: alive_out = 1;
            {6'd37, 6'd36}: alive_out = 1;
            {6'd37, 6'd37}: alive_out = 1;
            {6'd38, 6'd27}: alive_out = 1;
            {6'd38, 6'd30}: alive_out = 1;
            {6'd38, 6'd34}: alive_out = 1;
            {6'd38, 6'd37}: alive_out = 1;
            {6'd39, 6'd28}: alive_out = 1;
            {6'd39, 6'd29}: alive_out = 1;
            {6'd39, 6'd30}: alive_out = 1;
            {6'd39, 6'd34}: alive_out = 1;
            {6'd39, 6'd35}: alive_out = 1;
            {6'd39, 6'd36}: alive_out = 1;
            {6'd44, 6'd11}: alive_out = 1;
            {6'd44, 6'd12}: alive_out = 1;
            {6'd44, 6'd25}: alive_out = 1;
            {6'd44, 6'd26}: alive_out = 1;
            {6'd45, 6'd11}: alive_out = 1;
            {6'd45, 6'd12}: alive_out = 1;
            {6'd45, 6'd15}: alive_out = 1;
            {6'd45, 6'd16}: alive_out = 1;
            {6'd45, 6'd22}: alive_out = 1;
            {6'd45, 6'd23}: alive_out = 1;
            {6'd45, 6'd25}: alive_out = 1;
            {6'd45, 6'd26}: alive_out = 1;
            {6'd46, 6'd15}: alive_out = 1;
            {6'd46, 6'd16}: alive_out = 1;
            {6'd46, 6'd22}: alive_out = 1;
            {6'd46, 6'd23}: alive_out = 1;
            {6'd47, 6'd28}: alive_out = 1;
            {6'd47, 6'd29}: alive_out = 1;
            {6'd48, 6'd28}: alive_out = 1;
            {6'd48, 6'd29}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module simkinglidergun(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd14}: alive_out = 1;
            {6'd8, 6'd15}: alive_out = 1;
            {6'd9, 6'd14}: alive_out = 1;
            {6'd9, 6'd15}: alive_out = 1;
            {6'd12, 6'd16}: alive_out = 1;
            {6'd12, 6'd17}: alive_out = 1;
            {6'd13, 6'd16}: alive_out = 1;
            {6'd13, 6'd17}: alive_out = 1;
            {6'd15, 6'd14}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd16, 6'd14}: alive_out = 1;
            {6'd16, 6'd15}: alive_out = 1;
            {6'd28, 6'd23}: alive_out = 1;
            {6'd28, 6'd24}: alive_out = 1;
            {6'd29, 6'd19}: alive_out = 1;
            {6'd29, 6'd20}: alive_out = 1;
            {6'd29, 6'd21}: alive_out = 1;
            {6'd29, 6'd23}: alive_out = 1;
            {6'd29, 6'd25}: alive_out = 1;
            {6'd30, 6'd18}: alive_out = 1;
            {6'd30, 6'd21}: alive_out = 1;
            {6'd30, 6'd25}: alive_out = 1;
            {6'd31, 6'd18}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd25}: alive_out = 1;
            {6'd31, 6'd26}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd22}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd35, 6'd21}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd39, 6'd20}: alive_out = 1;
            {6'd39, 6'd21}: alive_out = 1;
            {6'd40, 6'd20}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module lobster(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd12, 6'd26}: alive_out = 1;
            {6'd12, 6'd32}: alive_out = 1;
            {6'd13, 6'd25}: alive_out = 1;
            {6'd13, 6'd31}: alive_out = 1;
            {6'd13, 6'd32}: alive_out = 1;
            {6'd14, 6'd25}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd15, 6'd26}: alive_out = 1;
            {6'd15, 6'd31}: alive_out = 1;
            {6'd16, 6'd26}: alive_out = 1;
            {6'd16, 6'd35}: alive_out = 1;
            {6'd16, 6'd36}: alive_out = 1;
            {6'd17, 6'd22}: alive_out = 1;
            {6'd17, 6'd23}: alive_out = 1;
            {6'd17, 6'd27}: alive_out = 1;
            {6'd17, 6'd33}: alive_out = 1;
            {6'd17, 6'd35}: alive_out = 1;
            {6'd18, 6'd21}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd29}: alive_out = 1;
            {6'd18, 6'd30}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd30}: alive_out = 1;
            {6'd19, 6'd34}: alive_out = 1;
            {6'd20, 6'd14}: alive_out = 1;
            {6'd20, 6'd15}: alive_out = 1;
            {6'd20, 6'd19}: alive_out = 1;
            {6'd20, 6'd21}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd27}: alive_out = 1;
            {6'd21, 6'd14}: alive_out = 1;
            {6'd21, 6'd15}: alive_out = 1;
            {6'd21, 6'd21}: alive_out = 1;
            {6'd21, 6'd28}: alive_out = 1;
            {6'd21, 6'd31}: alive_out = 1;
            {6'd22, 6'd18}: alive_out = 1;
            {6'd22, 6'd21}: alive_out = 1;
            {6'd22, 6'd28}: alive_out = 1;
            {6'd22, 6'd29}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd22, 6'd36}: alive_out = 1;
            {6'd23, 6'd12}: alive_out = 1;
            {6'd23, 6'd17}: alive_out = 1;
            {6'd23, 6'd19}: alive_out = 1;
            {6'd23, 6'd20}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd24, 6'd12}: alive_out = 1;
            {6'd24, 6'd14}: alive_out = 1;
            {6'd24, 6'd16}: alive_out = 1;
            {6'd24, 6'd17}: alive_out = 1;
            {6'd24, 6'd30}: alive_out = 1;
            {6'd25, 6'd12}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd25, 6'd16}: alive_out = 1;
            {6'd25, 6'd18}: alive_out = 1;
            {6'd25, 6'd31}: alive_out = 1;
            {6'd26, 6'd31}: alive_out = 1;
            {6'd27, 6'd26}: alive_out = 1;
            {6'd27, 6'd27}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd27, 6'd30}: alive_out = 1;
            {6'd28, 6'd25}: alive_out = 1;
            {6'd28, 6'd29}: alive_out = 1;
            {6'd29, 6'd25}: alive_out = 1;
            {6'd29, 6'd28}: alive_out = 1;
            {6'd31, 6'd23}: alive_out = 1;
            {6'd31, 6'd26}: alive_out = 1;
            {6'd32, 6'd24}: alive_out = 1;
            {6'd32, 6'd25}: alive_out = 1;
            {6'd33, 6'd23}: alive_out = 1;
            {6'd33, 6'd24}: alive_out = 1;
            {6'd34, 6'd27}: alive_out = 1;
            {6'd34, 6'd28}: alive_out = 1;
            {6'd35, 6'd24}: alive_out = 1;
            {6'd35, 6'd27}: alive_out = 1;
            {6'd35, 6'd28}: alive_out = 1;
            {6'd36, 6'd23}: alive_out = 1;
            {6'd37, 6'd23}: alive_out = 1;
            {6'd37, 6'd24}: alive_out = 1;
            {6'd37, 6'd25}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module snark(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd16, 6'd21}: alive_out = 1;
            {6'd17, 6'd21}: alive_out = 1;
            {6'd17, 6'd22}: alive_out = 1;
            {6'd17, 6'd23}: alive_out = 1;
            {6'd18, 6'd24}: alive_out = 1;
            {6'd18, 6'd27}: alive_out = 1;
            {6'd19, 6'd23}: alive_out = 1;
            {6'd19, 6'd24}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd27}: alive_out = 1;
            {6'd20, 6'd28}: alive_out = 1;
            {6'd22, 6'd13}: alive_out = 1;
            {6'd22, 6'd14}: alive_out = 1;
            {6'd22, 6'd16}: alive_out = 1;
            {6'd22, 6'd17}: alive_out = 1;
            {6'd23, 6'd13}: alive_out = 1;
            {6'd23, 6'd14}: alive_out = 1;
            {6'd23, 6'd16}: alive_out = 1;
            {6'd24, 6'd16}: alive_out = 1;
            {6'd25, 6'd16}: alive_out = 1;
            {6'd25, 6'd17}: alive_out = 1;
            {6'd25, 6'd18}: alive_out = 1;
            {6'd25, 6'd22}: alive_out = 1;
            {6'd25, 6'd23}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd15}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd23}: alive_out = 1;
            {6'd27, 6'd13}: alive_out = 1;
            {6'd27, 6'd16}: alive_out = 1;
            {6'd27, 6'd17}: alive_out = 1;
            {6'd27, 6'd18}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd28, 6'd13}: alive_out = 1;
            {6'd28, 6'd14}: alive_out = 1;
            {6'd28, 6'd16}: alive_out = 1;
            {6'd28, 6'd25}: alive_out = 1;
            {6'd28, 6'd26}: alive_out = 1;
            {6'd29, 6'd14}: alive_out = 1;
            {6'd29, 6'd17}: alive_out = 1;
            {6'd29, 6'd18}: alive_out = 1;
            {6'd29, 6'd19}: alive_out = 1;
            {6'd29, 6'd25}: alive_out = 1;
            {6'd29, 6'd27}: alive_out = 1;
            {6'd30, 6'd14}: alive_out = 1;
            {6'd30, 6'd20}: alive_out = 1;
            {6'd30, 6'd27}: alive_out = 1;
            {6'd31, 6'd15}: alive_out = 1;
            {6'd31, 6'd16}: alive_out = 1;
            {6'd31, 6'd17}: alive_out = 1;
            {6'd31, 6'd18}: alive_out = 1;
            {6'd31, 6'd19}: alive_out = 1;
            {6'd31, 6'd27}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd32, 6'd17}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module dinnertableextension(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd28}: alive_out = 1;
            {6'd9, 6'd17}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd9, 6'd26}: alive_out = 1;
            {6'd9, 6'd27}: alive_out = 1;
            {6'd9, 6'd28}: alive_out = 1;
            {6'd10, 6'd18}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd11, 6'd18}: alive_out = 1;
            {6'd11, 6'd20}: alive_out = 1;
            {6'd11, 6'd25}: alive_out = 1;
            {6'd11, 6'd26}: alive_out = 1;
            {6'd11, 6'd32}: alive_out = 1;
            {6'd12, 6'd19}: alive_out = 1;
            {6'd12, 6'd20}: alive_out = 1;
            {6'd12, 6'd30}: alive_out = 1;
            {6'd12, 6'd31}: alive_out = 1;
            {6'd12, 6'd32}: alive_out = 1;
            {6'd13, 6'd14}: alive_out = 1;
            {6'd13, 6'd15}: alive_out = 1;
            {6'd13, 6'd23}: alive_out = 1;
            {6'd13, 6'd24}: alive_out = 1;
            {6'd13, 6'd29}: alive_out = 1;
            {6'd14, 6'd15}: alive_out = 1;
            {6'd14, 6'd23}: alive_out = 1;
            {6'd14, 6'd24}: alive_out = 1;
            {6'd14, 6'd29}: alive_out = 1;
            {6'd14, 6'd30}: alive_out = 1;
            {6'd14, 6'd36}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd15, 6'd17}: alive_out = 1;
            {6'd15, 6'd23}: alive_out = 1;
            {6'd15, 6'd24}: alive_out = 1;
            {6'd15, 6'd34}: alive_out = 1;
            {6'd15, 6'd35}: alive_out = 1;
            {6'd15, 6'd36}: alive_out = 1;
            {6'd16, 6'd16}: alive_out = 1;
            {6'd16, 6'd17}: alive_out = 1;
            {6'd16, 6'd26}: alive_out = 1;
            {6'd16, 6'd27}: alive_out = 1;
            {6'd16, 6'd33}: alive_out = 1;
            {6'd17, 6'd11}: alive_out = 1;
            {6'd17, 6'd12}: alive_out = 1;
            {6'd17, 6'd19}: alive_out = 1;
            {6'd17, 6'd20}: alive_out = 1;
            {6'd17, 6'd26}: alive_out = 1;
            {6'd17, 6'd27}: alive_out = 1;
            {6'd17, 6'd33}: alive_out = 1;
            {6'd17, 6'd34}: alive_out = 1;
            {6'd17, 6'd40}: alive_out = 1;
            {6'd18, 6'd12}: alive_out = 1;
            {6'd18, 6'd19}: alive_out = 1;
            {6'd18, 6'd20}: alive_out = 1;
            {6'd18, 6'd26}: alive_out = 1;
            {6'd18, 6'd27}: alive_out = 1;
            {6'd18, 6'd38}: alive_out = 1;
            {6'd18, 6'd39}: alive_out = 1;
            {6'd18, 6'd40}: alive_out = 1;
            {6'd19, 6'd12}: alive_out = 1;
            {6'd19, 6'd14}: alive_out = 1;
            {6'd19, 6'd19}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd19, 6'd31}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd19, 6'd37}: alive_out = 1;
            {6'd20, 6'd13}: alive_out = 1;
            {6'd20, 6'd14}: alive_out = 1;
            {6'd20, 6'd24}: alive_out = 1;
            {6'd20, 6'd25}: alive_out = 1;
            {6'd20, 6'd31}: alive_out = 1;
            {6'd20, 6'd32}: alive_out = 1;
            {6'd20, 6'd37}: alive_out = 1;
            {6'd20, 6'd38}: alive_out = 1;
            {6'd21, 6'd8}: alive_out = 1;
            {6'd21, 6'd9}: alive_out = 1;
            {6'd21, 6'd17}: alive_out = 1;
            {6'd21, 6'd18}: alive_out = 1;
            {6'd21, 6'd24}: alive_out = 1;
            {6'd21, 6'd25}: alive_out = 1;
            {6'd21, 6'd31}: alive_out = 1;
            {6'd21, 6'd32}: alive_out = 1;
            {6'd22, 6'd9}: alive_out = 1;
            {6'd22, 6'd17}: alive_out = 1;
            {6'd22, 6'd18}: alive_out = 1;
            {6'd22, 6'd24}: alive_out = 1;
            {6'd22, 6'd25}: alive_out = 1;
            {6'd22, 6'd34}: alive_out = 1;
            {6'd22, 6'd35}: alive_out = 1;
            {6'd23, 6'd9}: alive_out = 1;
            {6'd23, 6'd11}: alive_out = 1;
            {6'd23, 6'd17}: alive_out = 1;
            {6'd23, 6'd18}: alive_out = 1;
            {6'd23, 6'd27}: alive_out = 1;
            {6'd23, 6'd28}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd24, 6'd10}: alive_out = 1;
            {6'd24, 6'd11}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd21}: alive_out = 1;
            {6'd24, 6'd27}: alive_out = 1;
            {6'd24, 6'd28}: alive_out = 1;
            {6'd24, 6'd34}: alive_out = 1;
            {6'd24, 6'd35}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd25, 6'd14}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd21}: alive_out = 1;
            {6'd25, 6'd27}: alive_out = 1;
            {6'd25, 6'd28}: alive_out = 1;
            {6'd25, 6'd38}: alive_out = 1;
            {6'd25, 6'd39}: alive_out = 1;
            {6'd26, 6'd13}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd21}: alive_out = 1;
            {6'd26, 6'd32}: alive_out = 1;
            {6'd26, 6'd33}: alive_out = 1;
            {6'd26, 6'd38}: alive_out = 1;
            {6'd26, 6'd40}: alive_out = 1;
            {6'd27, 6'd13}: alive_out = 1;
            {6'd27, 6'd14}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd27, 6'd26}: alive_out = 1;
            {6'd27, 6'd32}: alive_out = 1;
            {6'd27, 6'd33}: alive_out = 1;
            {6'd27, 6'd40}: alive_out = 1;
            {6'd28, 6'd18}: alive_out = 1;
            {6'd28, 6'd19}: alive_out = 1;
            {6'd28, 6'd25}: alive_out = 1;
            {6'd28, 6'd26}: alive_out = 1;
            {6'd28, 6'd32}: alive_out = 1;
            {6'd28, 6'd33}: alive_out = 1;
            {6'd28, 6'd40}: alive_out = 1;
            {6'd28, 6'd41}: alive_out = 1;
            {6'd29, 6'd11}: alive_out = 1;
            {6'd29, 6'd12}: alive_out = 1;
            {6'd29, 6'd18}: alive_out = 1;
            {6'd29, 6'd19}: alive_out = 1;
            {6'd29, 6'd25}: alive_out = 1;
            {6'd29, 6'd26}: alive_out = 1;
            {6'd29, 6'd35}: alive_out = 1;
            {6'd29, 6'd36}: alive_out = 1;
            {6'd30, 6'd12}: alive_out = 1;
            {6'd30, 6'd18}: alive_out = 1;
            {6'd30, 6'd19}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd29}: alive_out = 1;
            {6'd30, 6'd35}: alive_out = 1;
            {6'd30, 6'd37}: alive_out = 1;
            {6'd31, 6'd9}: alive_out = 1;
            {6'd31, 6'd10}: alive_out = 1;
            {6'd31, 6'd11}: alive_out = 1;
            {6'd31, 6'd21}: alive_out = 1;
            {6'd31, 6'd22}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd31, 6'd37}: alive_out = 1;
            {6'd32, 6'd9}: alive_out = 1;
            {6'd32, 6'd15}: alive_out = 1;
            {6'd32, 6'd16}: alive_out = 1;
            {6'd32, 6'd21}: alive_out = 1;
            {6'd32, 6'd22}: alive_out = 1;
            {6'd32, 6'd28}: alive_out = 1;
            {6'd32, 6'd29}: alive_out = 1;
            {6'd32, 6'd37}: alive_out = 1;
            {6'd32, 6'd38}: alive_out = 1;
            {6'd33, 6'd16}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd22}: alive_out = 1;
            {6'd33, 6'd32}: alive_out = 1;
            {6'd33, 6'd33}: alive_out = 1;
            {6'd34, 6'd13}: alive_out = 1;
            {6'd34, 6'd14}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd26}: alive_out = 1;
            {6'd34, 6'd27}: alive_out = 1;
            {6'd34, 6'd32}: alive_out = 1;
            {6'd34, 6'd34}: alive_out = 1;
            {6'd35, 6'd13}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd35, 6'd20}: alive_out = 1;
            {6'd35, 6'd26}: alive_out = 1;
            {6'd35, 6'd27}: alive_out = 1;
            {6'd35, 6'd34}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd36, 6'd26}: alive_out = 1;
            {6'd36, 6'd27}: alive_out = 1;
            {6'd36, 6'd34}: alive_out = 1;
            {6'd36, 6'd35}: alive_out = 1;
            {6'd37, 6'd17}: alive_out = 1;
            {6'd37, 6'd18}: alive_out = 1;
            {6'd37, 6'd19}: alive_out = 1;
            {6'd37, 6'd29}: alive_out = 1;
            {6'd37, 6'd30}: alive_out = 1;
            {6'd38, 6'd17}: alive_out = 1;
            {6'd38, 6'd23}: alive_out = 1;
            {6'd38, 6'd24}: alive_out = 1;
            {6'd38, 6'd29}: alive_out = 1;
            {6'd38, 6'd31}: alive_out = 1;
            {6'd39, 6'd24}: alive_out = 1;
            {6'd39, 6'd31}: alive_out = 1;
            {6'd40, 6'd21}: alive_out = 1;
            {6'd40, 6'd22}: alive_out = 1;
            {6'd40, 6'd23}: alive_out = 1;
            {6'd40, 6'd31}: alive_out = 1;
            {6'd40, 6'd32}: alive_out = 1;
            {6'd41, 6'd21}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module copperhead(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd21, 6'd22}: alive_out = 1;
            {6'd21, 6'd23}: alive_out = 1;
            {6'd21, 6'd24}: alive_out = 1;
            {6'd22, 6'd19}: alive_out = 1;
            {6'd22, 6'd25}: alive_out = 1;
            {6'd23, 6'd19}: alive_out = 1;
            {6'd23, 6'd22}: alive_out = 1;
            {6'd23, 6'd25}: alive_out = 1;
            {6'd23, 6'd26}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd21}: alive_out = 1;
            {6'd24, 6'd26}: alive_out = 1;
            {6'd24, 6'd27}: alive_out = 1;
            {6'd24, 6'd28}: alive_out = 1;
            {6'd25, 6'd20}: alive_out = 1;
            {6'd25, 6'd21}: alive_out = 1;
            {6'd25, 6'd26}: alive_out = 1;
            {6'd25, 6'd27}: alive_out = 1;
            {6'd25, 6'd28}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd22}: alive_out = 1;
            {6'd26, 6'd25}: alive_out = 1;
            {6'd26, 6'd26}: alive_out = 1;
            {6'd27, 6'd19}: alive_out = 1;
            {6'd27, 6'd25}: alive_out = 1;
            {6'd28, 6'd22}: alive_out = 1;
            {6'd28, 6'd23}: alive_out = 1;
            {6'd28, 6'd24}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module p50glidershuttle(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd8, 6'd24}: alive_out = 1;
            {6'd9, 6'd23}: alive_out = 1;
            {6'd9, 6'd25}: alive_out = 1;
            {6'd10, 6'd18}: alive_out = 1;
            {6'd10, 6'd23}: alive_out = 1;
            {6'd10, 6'd25}: alive_out = 1;
            {6'd11, 6'd17}: alive_out = 1;
            {6'd11, 6'd19}: alive_out = 1;
            {6'd11, 6'd22}: alive_out = 1;
            {6'd11, 6'd23}: alive_out = 1;
            {6'd11, 6'd25}: alive_out = 1;
            {6'd11, 6'd26}: alive_out = 1;
            {6'd11, 6'd29}: alive_out = 1;
            {6'd11, 6'd30}: alive_out = 1;
            {6'd12, 6'd18}: alive_out = 1;
            {6'd12, 6'd22}: alive_out = 1;
            {6'd12, 6'd28}: alive_out = 1;
            {6'd12, 6'd31}: alive_out = 1;
            {6'd13, 6'd23}: alive_out = 1;
            {6'd13, 6'd24}: alive_out = 1;
            {6'd13, 6'd25}: alive_out = 1;
            {6'd13, 6'd30}: alive_out = 1;
            {6'd13, 6'd33}: alive_out = 1;
            {6'd14, 6'd16}: alive_out = 1;
            {6'd14, 6'd17}: alive_out = 1;
            {6'd14, 6'd18}: alive_out = 1;
            {6'd14, 6'd19}: alive_out = 1;
            {6'd14, 6'd20}: alive_out = 1;
            {6'd14, 6'd25}: alive_out = 1;
            {6'd14, 6'd28}: alive_out = 1;
            {6'd14, 6'd30}: alive_out = 1;
            {6'd14, 6'd32}: alive_out = 1;
            {6'd14, 6'd33}: alive_out = 1;
            {6'd15, 6'd15}: alive_out = 1;
            {6'd15, 6'd20}: alive_out = 1;
            {6'd15, 6'd26}: alive_out = 1;
            {6'd15, 6'd27}: alive_out = 1;
            {6'd15, 6'd30}: alive_out = 1;
            {6'd15, 6'd34}: alive_out = 1;
            {6'd15, 6'd35}: alive_out = 1;
            {6'd16, 6'd14}: alive_out = 1;
            {6'd16, 6'd17}: alive_out = 1;
            {6'd16, 6'd29}: alive_out = 1;
            {6'd16, 6'd30}: alive_out = 1;
            {6'd16, 6'd34}: alive_out = 1;
            {6'd17, 6'd11}: alive_out = 1;
            {6'd17, 6'd14}: alive_out = 1;
            {6'd17, 6'd16}: alive_out = 1;
            {6'd17, 6'd17}: alive_out = 1;
            {6'd17, 6'd36}: alive_out = 1;
            {6'd18, 6'd10}: alive_out = 1;
            {6'd18, 6'd12}: alive_out = 1;
            {6'd18, 6'd14}: alive_out = 1;
            {6'd18, 6'd20}: alive_out = 1;
            {6'd18, 6'd32}: alive_out = 1;
            {6'd18, 6'd33}: alive_out = 1;
            {6'd18, 6'd34}: alive_out = 1;
            {6'd18, 6'd35}: alive_out = 1;
            {6'd18, 6'd37}: alive_out = 1;
            {6'd19, 6'd11}: alive_out = 1;
            {6'd19, 6'd14}: alive_out = 1;
            {6'd19, 6'd19}: alive_out = 1;
            {6'd19, 6'd21}: alive_out = 1;
            {6'd19, 6'd26}: alive_out = 1;
            {6'd19, 6'd32}: alive_out = 1;
            {6'd19, 6'd37}: alive_out = 1;
            {6'd20, 6'd14}: alive_out = 1;
            {6'd20, 6'd15}: alive_out = 1;
            {6'd20, 6'd18}: alive_out = 1;
            {6'd20, 6'd21}: alive_out = 1;
            {6'd20, 6'd24}: alive_out = 1;
            {6'd20, 6'd26}: alive_out = 1;
            {6'd20, 6'd34}: alive_out = 1;
            {6'd20, 6'd36}: alive_out = 1;
            {6'd21, 6'd19}: alive_out = 1;
            {6'd21, 6'd20}: alive_out = 1;
            {6'd21, 6'd25}: alive_out = 1;
            {6'd21, 6'd26}: alive_out = 1;
            {6'd21, 6'd33}: alive_out = 1;
            {6'd22, 6'd11}: alive_out = 1;
            {6'd22, 6'd12}: alive_out = 1;
            {6'd22, 6'd33}: alive_out = 1;
            {6'd22, 6'd37}: alive_out = 1;
            {6'd23, 6'd9}: alive_out = 1;
            {6'd23, 6'd10}: alive_out = 1;
            {6'd23, 6'd11}: alive_out = 1;
            {6'd23, 6'd13}: alive_out = 1;
            {6'd23, 6'd34}: alive_out = 1;
            {6'd23, 6'd35}: alive_out = 1;
            {6'd23, 6'd37}: alive_out = 1;
            {6'd23, 6'd38}: alive_out = 1;
            {6'd23, 6'd39}: alive_out = 1;
            {6'd24, 6'd8}: alive_out = 1;
            {6'd24, 6'd13}: alive_out = 1;
            {6'd24, 6'd20}: alive_out = 1;
            {6'd24, 6'd35}: alive_out = 1;
            {6'd24, 6'd40}: alive_out = 1;
            {6'd25, 6'd9}: alive_out = 1;
            {6'd25, 6'd10}: alive_out = 1;
            {6'd25, 6'd11}: alive_out = 1;
            {6'd25, 6'd13}: alive_out = 1;
            {6'd25, 6'd14}: alive_out = 1;
            {6'd25, 6'd21}: alive_out = 1;
            {6'd25, 6'd35}: alive_out = 1;
            {6'd25, 6'd37}: alive_out = 1;
            {6'd25, 6'd38}: alive_out = 1;
            {6'd25, 6'd39}: alive_out = 1;
            {6'd26, 6'd11}: alive_out = 1;
            {6'd26, 6'd15}: alive_out = 1;
            {6'd26, 6'd19}: alive_out = 1;
            {6'd26, 6'd20}: alive_out = 1;
            {6'd26, 6'd21}: alive_out = 1;
            {6'd26, 6'd36}: alive_out = 1;
            {6'd26, 6'd37}: alive_out = 1;
            {6'd27, 6'd15}: alive_out = 1;
            {6'd27, 6'd28}: alive_out = 1;
            {6'd27, 6'd29}: alive_out = 1;
            {6'd28, 6'd12}: alive_out = 1;
            {6'd28, 6'd14}: alive_out = 1;
            {6'd28, 6'd27}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd28, 6'd33}: alive_out = 1;
            {6'd28, 6'd34}: alive_out = 1;
            {6'd29, 6'd11}: alive_out = 1;
            {6'd29, 6'd16}: alive_out = 1;
            {6'd29, 6'd27}: alive_out = 1;
            {6'd29, 6'd29}: alive_out = 1;
            {6'd29, 6'd34}: alive_out = 1;
            {6'd29, 6'd37}: alive_out = 1;
            {6'd30, 6'd11}: alive_out = 1;
            {6'd30, 6'd13}: alive_out = 1;
            {6'd30, 6'd14}: alive_out = 1;
            {6'd30, 6'd15}: alive_out = 1;
            {6'd30, 6'd16}: alive_out = 1;
            {6'd30, 6'd28}: alive_out = 1;
            {6'd30, 6'd34}: alive_out = 1;
            {6'd30, 6'd36}: alive_out = 1;
            {6'd30, 6'd38}: alive_out = 1;
            {6'd31, 6'd12}: alive_out = 1;
            {6'd31, 6'd31}: alive_out = 1;
            {6'd31, 6'd32}: alive_out = 1;
            {6'd31, 6'd34}: alive_out = 1;
            {6'd31, 6'd37}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd18}: alive_out = 1;
            {6'd32, 6'd19}: alive_out = 1;
            {6'd32, 6'd31}: alive_out = 1;
            {6'd32, 6'd34}: alive_out = 1;
            {6'd33, 6'd13}: alive_out = 1;
            {6'd33, 6'd14}: alive_out = 1;
            {6'd33, 6'd18}: alive_out = 1;
            {6'd33, 6'd21}: alive_out = 1;
            {6'd33, 6'd22}: alive_out = 1;
            {6'd33, 6'd28}: alive_out = 1;
            {6'd33, 6'd33}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd16}: alive_out = 1;
            {6'd34, 6'd18}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd34, 6'd23}: alive_out = 1;
            {6'd34, 6'd28}: alive_out = 1;
            {6'd34, 6'd29}: alive_out = 1;
            {6'd34, 6'd30}: alive_out = 1;
            {6'd34, 6'd31}: alive_out = 1;
            {6'd34, 6'd32}: alive_out = 1;
            {6'd35, 6'd15}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd23}: alive_out = 1;
            {6'd35, 6'd24}: alive_out = 1;
            {6'd35, 6'd25}: alive_out = 1;
            {6'd36, 6'd17}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd36, 6'd26}: alive_out = 1;
            {6'd36, 6'd30}: alive_out = 1;
            {6'd37, 6'd18}: alive_out = 1;
            {6'd37, 6'd19}: alive_out = 1;
            {6'd37, 6'd22}: alive_out = 1;
            {6'd37, 6'd23}: alive_out = 1;
            {6'd37, 6'd25}: alive_out = 1;
            {6'd37, 6'd26}: alive_out = 1;
            {6'd37, 6'd29}: alive_out = 1;
            {6'd37, 6'd31}: alive_out = 1;
            {6'd38, 6'd23}: alive_out = 1;
            {6'd38, 6'd25}: alive_out = 1;
            {6'd38, 6'd30}: alive_out = 1;
            {6'd39, 6'd23}: alive_out = 1;
            {6'd39, 6'd25}: alive_out = 1;
            {6'd40, 6'd24}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module hectic(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd5, 6'd10}: alive_out = 1;
            {6'd5, 6'd11}: alive_out = 1;
            {6'd6, 6'd10}: alive_out = 1;
            {6'd6, 6'd11}: alive_out = 1;
            {6'd10, 6'd10}: alive_out = 1;
            {6'd11, 6'd9}: alive_out = 1;
            {6'd11, 6'd11}: alive_out = 1;
            {6'd12, 6'd8}: alive_out = 1;
            {6'd12, 6'd12}: alive_out = 1;
            {6'd13, 6'd9}: alive_out = 1;
            {6'd13, 6'd10}: alive_out = 1;
            {6'd13, 6'd11}: alive_out = 1;
            {6'd14, 6'd7}: alive_out = 1;
            {6'd14, 6'd8}: alive_out = 1;
            {6'd14, 6'd12}: alive_out = 1;
            {6'd14, 6'd13}: alive_out = 1;
            {6'd17, 6'd21}: alive_out = 1;
            {6'd18, 6'd19}: alive_out = 1;
            {6'd18, 6'd21}: alive_out = 1;
            {6'd19, 6'd18}: alive_out = 1;
            {6'd19, 6'd20}: alive_out = 1;
            {6'd20, 6'd17}: alive_out = 1;
            {6'd20, 6'd20}: alive_out = 1;
            {6'd20, 6'd22}: alive_out = 1;
            {6'd20, 6'd23}: alive_out = 1;
            {6'd21, 6'd12}: alive_out = 1;
            {6'd21, 6'd13}: alive_out = 1;
            {6'd21, 6'd18}: alive_out = 1;
            {6'd21, 6'd20}: alive_out = 1;
            {6'd21, 6'd22}: alive_out = 1;
            {6'd21, 6'd23}: alive_out = 1;
            {6'd22, 6'd13}: alive_out = 1;
            {6'd22, 6'd14}: alive_out = 1;
            {6'd22, 6'd19}: alive_out = 1;
            {6'd22, 6'd21}: alive_out = 1;
            {6'd23, 6'd12}: alive_out = 1;
            {6'd23, 6'd21}: alive_out = 1;
            {6'd25, 6'd7}: alive_out = 1;
            {6'd25, 6'd16}: alive_out = 1;
            {6'd26, 6'd7}: alive_out = 1;
            {6'd26, 6'd9}: alive_out = 1;
            {6'd26, 6'd14}: alive_out = 1;
            {6'd26, 6'd15}: alive_out = 1;
            {6'd27, 6'd5}: alive_out = 1;
            {6'd27, 6'd6}: alive_out = 1;
            {6'd27, 6'd8}: alive_out = 1;
            {6'd27, 6'd10}: alive_out = 1;
            {6'd27, 6'd15}: alive_out = 1;
            {6'd27, 6'd16}: alive_out = 1;
            {6'd28, 6'd5}: alive_out = 1;
            {6'd28, 6'd6}: alive_out = 1;
            {6'd28, 6'd8}: alive_out = 1;
            {6'd28, 6'd11}: alive_out = 1;
            {6'd29, 6'd8}: alive_out = 1;
            {6'd29, 6'd10}: alive_out = 1;
            {6'd30, 6'd7}: alive_out = 1;
            {6'd30, 6'd9}: alive_out = 1;
            {6'd31, 6'd7}: alive_out = 1;
            {6'd34, 6'd15}: alive_out = 1;
            {6'd34, 6'd16}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd34, 6'd21}: alive_out = 1;
            {6'd35, 6'd17}: alive_out = 1;
            {6'd35, 6'd18}: alive_out = 1;
            {6'd35, 6'd19}: alive_out = 1;
            {6'd36, 6'd16}: alive_out = 1;
            {6'd36, 6'd20}: alive_out = 1;
            {6'd37, 6'd17}: alive_out = 1;
            {6'd37, 6'd19}: alive_out = 1;
            {6'd38, 6'd18}: alive_out = 1;
            {6'd42, 6'd17}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd43, 6'd17}: alive_out = 1;
            {6'd43, 6'd18}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module p45engine(input wire[5:0] x_in,
               input wire[5:0] y_in,
               output logic alive_out);
    always_comb begin
        case ({x_in, y_in})
            {6'd4, 6'd19}: alive_out = 1;
            {6'd4, 6'd20}: alive_out = 1;
            {6'd5, 6'd20}: alive_out = 1;
            {6'd6, 6'd20}: alive_out = 1;
            {6'd6, 6'd22}: alive_out = 1;
            {6'd6, 6'd23}: alive_out = 1;
            {6'd7, 6'd15}: alive_out = 1;
            {6'd7, 6'd16}: alive_out = 1;
            {6'd7, 6'd21}: alive_out = 1;
            {6'd7, 6'd23}: alive_out = 1;
            {6'd8, 6'd16}: alive_out = 1;
            {6'd9, 6'd16}: alive_out = 1;
            {6'd9, 6'd18}: alive_out = 1;
            {6'd10, 6'd17}: alive_out = 1;
            {6'd10, 6'd18}: alive_out = 1;
            {6'd15, 6'd21}: alive_out = 1;
            {6'd15, 6'd24}: alive_out = 1;
            {6'd16, 6'd21}: alive_out = 1;
            {6'd16, 6'd24}: alive_out = 1;
            {6'd16, 6'd27}: alive_out = 1;
            {6'd16, 6'd28}: alive_out = 1;
            {6'd17, 6'd12}: alive_out = 1;
            {6'd17, 6'd13}: alive_out = 1;
            {6'd17, 6'd21}: alive_out = 1;
            {6'd17, 6'd24}: alive_out = 1;
            {6'd17, 6'd27}: alive_out = 1;
            {6'd17, 6'd28}: alive_out = 1;
            {6'd18, 6'd12}: alive_out = 1;
            {6'd18, 6'd13}: alive_out = 1;
            {6'd19, 6'd34}: alive_out = 1;
            {6'd20, 6'd32}: alive_out = 1;
            {6'd20, 6'd33}: alive_out = 1;
            {6'd20, 6'd34}: alive_out = 1;
            {6'd21, 6'd11}: alive_out = 1;
            {6'd21, 6'd12}: alive_out = 1;
            {6'd21, 6'd13}: alive_out = 1;
            {6'd21, 6'd31}: alive_out = 1;
            {6'd22, 6'd6}: alive_out = 1;
            {6'd22, 6'd7}: alive_out = 1;
            {6'd22, 6'd31}: alive_out = 1;
            {6'd22, 6'd32}: alive_out = 1;
            {6'd23, 6'd6}: alive_out = 1;
            {6'd23, 6'd37}: alive_out = 1;
            {6'd24, 6'd7}: alive_out = 1;
            {6'd24, 6'd11}: alive_out = 1;
            {6'd24, 6'd12}: alive_out = 1;
            {6'd24, 6'd13}: alive_out = 1;
            {6'd24, 6'd35}: alive_out = 1;
            {6'd24, 6'd36}: alive_out = 1;
            {6'd24, 6'd37}: alive_out = 1;
            {6'd25, 6'd4}: alive_out = 1;
            {6'd25, 6'd5}: alive_out = 1;
            {6'd25, 6'd6}: alive_out = 1;
            {6'd25, 6'd28}: alive_out = 1;
            {6'd25, 6'd29}: alive_out = 1;
            {6'd25, 6'd30}: alive_out = 1;
            {6'd25, 6'd34}: alive_out = 1;
            {6'd26, 6'd4}: alive_out = 1;
            {6'd26, 6'd35}: alive_out = 1;
            {6'd27, 6'd9}: alive_out = 1;
            {6'd27, 6'd10}: alive_out = 1;
            {6'd27, 6'd34}: alive_out = 1;
            {6'd27, 6'd35}: alive_out = 1;
            {6'd28, 6'd10}: alive_out = 1;
            {6'd28, 6'd28}: alive_out = 1;
            {6'd28, 6'd29}: alive_out = 1;
            {6'd28, 6'd30}: alive_out = 1;
            {6'd29, 6'd7}: alive_out = 1;
            {6'd29, 6'd8}: alive_out = 1;
            {6'd29, 6'd9}: alive_out = 1;
            {6'd30, 6'd7}: alive_out = 1;
            {6'd31, 6'd28}: alive_out = 1;
            {6'd31, 6'd29}: alive_out = 1;
            {6'd32, 6'd13}: alive_out = 1;
            {6'd32, 6'd14}: alive_out = 1;
            {6'd32, 6'd17}: alive_out = 1;
            {6'd32, 6'd20}: alive_out = 1;
            {6'd32, 6'd28}: alive_out = 1;
            {6'd32, 6'd29}: alive_out = 1;
            {6'd33, 6'd13}: alive_out = 1;
            {6'd33, 6'd14}: alive_out = 1;
            {6'd33, 6'd17}: alive_out = 1;
            {6'd33, 6'd20}: alive_out = 1;
            {6'd34, 6'd17}: alive_out = 1;
            {6'd34, 6'd20}: alive_out = 1;
            {6'd39, 6'd23}: alive_out = 1;
            {6'd39, 6'd24}: alive_out = 1;
            {6'd40, 6'd23}: alive_out = 1;
            {6'd40, 6'd25}: alive_out = 1;
            {6'd41, 6'd25}: alive_out = 1;
            {6'd42, 6'd18}: alive_out = 1;
            {6'd42, 6'd20}: alive_out = 1;
            {6'd42, 6'd25}: alive_out = 1;
            {6'd42, 6'd26}: alive_out = 1;
            {6'd43, 6'd18}: alive_out = 1;
            {6'd43, 6'd19}: alive_out = 1;
            {6'd43, 6'd21}: alive_out = 1;
            {6'd44, 6'd21}: alive_out = 1;
            {6'd45, 6'd21}: alive_out = 1;
            {6'd45, 6'd22}: alive_out = 1;

            default: alive_out = 0;
        endcase
    end
endmodule
`default_nettype wire
`default_nettype none
module seed_select(input wire[4:0] seed_idx,
                   input wire[5:0] x_in,
                   input wire[5:0] y_in,
                   output logic alive_out);
    logic alive[0:23];
    b52bomber s0(.x_in(x_in), .y_in(y_in), .alive_out(alive[0]));
    shipinabottle s1(.x_in(x_in), .y_in(y_in), .alive_out(alive[1]));
    loaflipflop s2(.x_in(x_in), .y_in(y_in), .alive_out(alive[2]));
    ringoffire s3(.x_in(x_in), .y_in(y_in), .alive_out(alive[3]));
    frothingpuffer s4(.x_in(x_in), .y_in(y_in), .alive_out(alive[4]));
    venetial_blinds s5(.x_in(x_in), .y_in(y_in), .alive_out(alive[5]));
    trafficcircle s6(.x_in(x_in), .y_in(y_in), .alive_out(alive[6]));
    superfountain s7(.x_in(x_in), .y_in(y_in), .alive_out(alive[7]));
    harvester s8(.x_in(x_in), .y_in(y_in), .alive_out(alive[8]));
    wickstrecher s9(.x_in(x_in), .y_in(y_in), .alive_out(alive[9]));
    rectifier s10(.x_in(x_in), .y_in(y_in), .alive_out(alive[10]));
    fly s11(.x_in(x_in), .y_in(y_in), .alive_out(alive[11]));
    spacefiller s12(.x_in(x_in), .y_in(y_in), .alive_out(alive[12]));
    pulsar s13(.x_in(x_in), .y_in(y_in), .alive_out(alive[13]));
    10cellinfinitegrowth s14(.x_in(x_in), .y_in(y_in), .alive_out(alive[14]));
    vacuumgun s15(.x_in(x_in), .y_in(y_in), .alive_out(alive[15]));
    simkinglidergun s16(.x_in(x_in), .y_in(y_in), .alive_out(alive[16]));
    lobster s17(.x_in(x_in), .y_in(y_in), .alive_out(alive[17]));
    snark s18(.x_in(x_in), .y_in(y_in), .alive_out(alive[18]));
    dinnertableextension s19(.x_in(x_in), .y_in(y_in), .alive_out(alive[19]));
    copperhead s20(.x_in(x_in), .y_in(y_in), .alive_out(alive[20]));
    p50glidershuttle s21(.x_in(x_in), .y_in(y_in), .alive_out(alive[21]));
    hectic s22(.x_in(x_in), .y_in(y_in), .alive_out(alive[22]));
    p45engine s23(.x_in(x_in), .y_in(y_in), .alive_out(alive[23]));
    assign alive_out = alive[seed_idx];
endmodule
`default_nettype wire
