`timescale 1ns / 1ps

module audio(input wire clk_100mhz,
             input wire rst_in,
             input wire miso_in,
             output logic cs_out, mosi_out, sclk_out);
endmodule

